magic
tech sky130A
magscale 1 2
timestamp 1697034114
<< pwell >>
rect -3521 -410 3521 410
<< nmos >>
rect -3325 -200 -3125 200
rect -3067 -200 -2867 200
rect -2809 -200 -2609 200
rect -2551 -200 -2351 200
rect -2293 -200 -2093 200
rect -2035 -200 -1835 200
rect -1777 -200 -1577 200
rect -1519 -200 -1319 200
rect -1261 -200 -1061 200
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
rect 1061 -200 1261 200
rect 1319 -200 1519 200
rect 1577 -200 1777 200
rect 1835 -200 2035 200
rect 2093 -200 2293 200
rect 2351 -200 2551 200
rect 2609 -200 2809 200
rect 2867 -200 3067 200
rect 3125 -200 3325 200
<< ndiff >>
rect -3383 188 -3325 200
rect -3383 -188 -3371 188
rect -3337 -188 -3325 188
rect -3383 -200 -3325 -188
rect -3125 188 -3067 200
rect -3125 -188 -3113 188
rect -3079 -188 -3067 188
rect -3125 -200 -3067 -188
rect -2867 188 -2809 200
rect -2867 -188 -2855 188
rect -2821 -188 -2809 188
rect -2867 -200 -2809 -188
rect -2609 188 -2551 200
rect -2609 -188 -2597 188
rect -2563 -188 -2551 188
rect -2609 -200 -2551 -188
rect -2351 188 -2293 200
rect -2351 -188 -2339 188
rect -2305 -188 -2293 188
rect -2351 -200 -2293 -188
rect -2093 188 -2035 200
rect -2093 -188 -2081 188
rect -2047 -188 -2035 188
rect -2093 -200 -2035 -188
rect -1835 188 -1777 200
rect -1835 -188 -1823 188
rect -1789 -188 -1777 188
rect -1835 -200 -1777 -188
rect -1577 188 -1519 200
rect -1577 -188 -1565 188
rect -1531 -188 -1519 188
rect -1577 -200 -1519 -188
rect -1319 188 -1261 200
rect -1319 -188 -1307 188
rect -1273 -188 -1261 188
rect -1319 -200 -1261 -188
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
rect 1261 188 1319 200
rect 1261 -188 1273 188
rect 1307 -188 1319 188
rect 1261 -200 1319 -188
rect 1519 188 1577 200
rect 1519 -188 1531 188
rect 1565 -188 1577 188
rect 1519 -200 1577 -188
rect 1777 188 1835 200
rect 1777 -188 1789 188
rect 1823 -188 1835 188
rect 1777 -200 1835 -188
rect 2035 188 2093 200
rect 2035 -188 2047 188
rect 2081 -188 2093 188
rect 2035 -200 2093 -188
rect 2293 188 2351 200
rect 2293 -188 2305 188
rect 2339 -188 2351 188
rect 2293 -200 2351 -188
rect 2551 188 2609 200
rect 2551 -188 2563 188
rect 2597 -188 2609 188
rect 2551 -200 2609 -188
rect 2809 188 2867 200
rect 2809 -188 2821 188
rect 2855 -188 2867 188
rect 2809 -200 2867 -188
rect 3067 188 3125 200
rect 3067 -188 3079 188
rect 3113 -188 3125 188
rect 3067 -200 3125 -188
rect 3325 188 3383 200
rect 3325 -188 3337 188
rect 3371 -188 3383 188
rect 3325 -200 3383 -188
<< ndiffc >>
rect -3371 -188 -3337 188
rect -3113 -188 -3079 188
rect -2855 -188 -2821 188
rect -2597 -188 -2563 188
rect -2339 -188 -2305 188
rect -2081 -188 -2047 188
rect -1823 -188 -1789 188
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect 1789 -188 1823 188
rect 2047 -188 2081 188
rect 2305 -188 2339 188
rect 2563 -188 2597 188
rect 2821 -188 2855 188
rect 3079 -188 3113 188
rect 3337 -188 3371 188
<< psubdiff >>
rect -3485 340 -3389 374
rect 3389 340 3485 374
rect -3485 278 -3451 340
rect 3451 278 3485 340
rect -3485 -340 -3451 -278
rect 3451 -340 3485 -278
rect -3485 -374 -3389 -340
rect 3389 -374 3485 -340
<< psubdiffcont >>
rect -3389 340 3389 374
rect -3485 -278 -3451 278
rect 3451 -278 3485 278
rect -3389 -374 3389 -340
<< poly >>
rect -3325 272 -3125 288
rect -3325 238 -3309 272
rect -3141 238 -3125 272
rect -3325 200 -3125 238
rect -3067 272 -2867 288
rect -3067 238 -3051 272
rect -2883 238 -2867 272
rect -3067 200 -2867 238
rect -2809 272 -2609 288
rect -2809 238 -2793 272
rect -2625 238 -2609 272
rect -2809 200 -2609 238
rect -2551 272 -2351 288
rect -2551 238 -2535 272
rect -2367 238 -2351 272
rect -2551 200 -2351 238
rect -2293 272 -2093 288
rect -2293 238 -2277 272
rect -2109 238 -2093 272
rect -2293 200 -2093 238
rect -2035 272 -1835 288
rect -2035 238 -2019 272
rect -1851 238 -1835 272
rect -2035 200 -1835 238
rect -1777 272 -1577 288
rect -1777 238 -1761 272
rect -1593 238 -1577 272
rect -1777 200 -1577 238
rect -1519 272 -1319 288
rect -1519 238 -1503 272
rect -1335 238 -1319 272
rect -1519 200 -1319 238
rect -1261 272 -1061 288
rect -1261 238 -1245 272
rect -1077 238 -1061 272
rect -1261 200 -1061 238
rect -1003 272 -803 288
rect -1003 238 -987 272
rect -819 238 -803 272
rect -1003 200 -803 238
rect -745 272 -545 288
rect -745 238 -729 272
rect -561 238 -545 272
rect -745 200 -545 238
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect 545 272 745 288
rect 545 238 561 272
rect 729 238 745 272
rect 545 200 745 238
rect 803 272 1003 288
rect 803 238 819 272
rect 987 238 1003 272
rect 803 200 1003 238
rect 1061 272 1261 288
rect 1061 238 1077 272
rect 1245 238 1261 272
rect 1061 200 1261 238
rect 1319 272 1519 288
rect 1319 238 1335 272
rect 1503 238 1519 272
rect 1319 200 1519 238
rect 1577 272 1777 288
rect 1577 238 1593 272
rect 1761 238 1777 272
rect 1577 200 1777 238
rect 1835 272 2035 288
rect 1835 238 1851 272
rect 2019 238 2035 272
rect 1835 200 2035 238
rect 2093 272 2293 288
rect 2093 238 2109 272
rect 2277 238 2293 272
rect 2093 200 2293 238
rect 2351 272 2551 288
rect 2351 238 2367 272
rect 2535 238 2551 272
rect 2351 200 2551 238
rect 2609 272 2809 288
rect 2609 238 2625 272
rect 2793 238 2809 272
rect 2609 200 2809 238
rect 2867 272 3067 288
rect 2867 238 2883 272
rect 3051 238 3067 272
rect 2867 200 3067 238
rect 3125 272 3325 288
rect 3125 238 3141 272
rect 3309 238 3325 272
rect 3125 200 3325 238
rect -3325 -238 -3125 -200
rect -3325 -272 -3309 -238
rect -3141 -272 -3125 -238
rect -3325 -288 -3125 -272
rect -3067 -238 -2867 -200
rect -3067 -272 -3051 -238
rect -2883 -272 -2867 -238
rect -3067 -288 -2867 -272
rect -2809 -238 -2609 -200
rect -2809 -272 -2793 -238
rect -2625 -272 -2609 -238
rect -2809 -288 -2609 -272
rect -2551 -238 -2351 -200
rect -2551 -272 -2535 -238
rect -2367 -272 -2351 -238
rect -2551 -288 -2351 -272
rect -2293 -238 -2093 -200
rect -2293 -272 -2277 -238
rect -2109 -272 -2093 -238
rect -2293 -288 -2093 -272
rect -2035 -238 -1835 -200
rect -2035 -272 -2019 -238
rect -1851 -272 -1835 -238
rect -2035 -288 -1835 -272
rect -1777 -238 -1577 -200
rect -1777 -272 -1761 -238
rect -1593 -272 -1577 -238
rect -1777 -288 -1577 -272
rect -1519 -238 -1319 -200
rect -1519 -272 -1503 -238
rect -1335 -272 -1319 -238
rect -1519 -288 -1319 -272
rect -1261 -238 -1061 -200
rect -1261 -272 -1245 -238
rect -1077 -272 -1061 -238
rect -1261 -288 -1061 -272
rect -1003 -238 -803 -200
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -1003 -288 -803 -272
rect -745 -238 -545 -200
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -745 -288 -545 -272
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
rect 545 -238 745 -200
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 545 -288 745 -272
rect 803 -238 1003 -200
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect 803 -288 1003 -272
rect 1061 -238 1261 -200
rect 1061 -272 1077 -238
rect 1245 -272 1261 -238
rect 1061 -288 1261 -272
rect 1319 -238 1519 -200
rect 1319 -272 1335 -238
rect 1503 -272 1519 -238
rect 1319 -288 1519 -272
rect 1577 -238 1777 -200
rect 1577 -272 1593 -238
rect 1761 -272 1777 -238
rect 1577 -288 1777 -272
rect 1835 -238 2035 -200
rect 1835 -272 1851 -238
rect 2019 -272 2035 -238
rect 1835 -288 2035 -272
rect 2093 -238 2293 -200
rect 2093 -272 2109 -238
rect 2277 -272 2293 -238
rect 2093 -288 2293 -272
rect 2351 -238 2551 -200
rect 2351 -272 2367 -238
rect 2535 -272 2551 -238
rect 2351 -288 2551 -272
rect 2609 -238 2809 -200
rect 2609 -272 2625 -238
rect 2793 -272 2809 -238
rect 2609 -288 2809 -272
rect 2867 -238 3067 -200
rect 2867 -272 2883 -238
rect 3051 -272 3067 -238
rect 2867 -288 3067 -272
rect 3125 -238 3325 -200
rect 3125 -272 3141 -238
rect 3309 -272 3325 -238
rect 3125 -288 3325 -272
<< polycont >>
rect -3309 238 -3141 272
rect -3051 238 -2883 272
rect -2793 238 -2625 272
rect -2535 238 -2367 272
rect -2277 238 -2109 272
rect -2019 238 -1851 272
rect -1761 238 -1593 272
rect -1503 238 -1335 272
rect -1245 238 -1077 272
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect 1077 238 1245 272
rect 1335 238 1503 272
rect 1593 238 1761 272
rect 1851 238 2019 272
rect 2109 238 2277 272
rect 2367 238 2535 272
rect 2625 238 2793 272
rect 2883 238 3051 272
rect 3141 238 3309 272
rect -3309 -272 -3141 -238
rect -3051 -272 -2883 -238
rect -2793 -272 -2625 -238
rect -2535 -272 -2367 -238
rect -2277 -272 -2109 -238
rect -2019 -272 -1851 -238
rect -1761 -272 -1593 -238
rect -1503 -272 -1335 -238
rect -1245 -272 -1077 -238
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
rect 1077 -272 1245 -238
rect 1335 -272 1503 -238
rect 1593 -272 1761 -238
rect 1851 -272 2019 -238
rect 2109 -272 2277 -238
rect 2367 -272 2535 -238
rect 2625 -272 2793 -238
rect 2883 -272 3051 -238
rect 3141 -272 3309 -238
<< locali >>
rect -3485 340 -3389 374
rect 3389 340 3485 374
rect -3485 278 -3451 340
rect 3451 278 3485 340
rect -3325 238 -3309 272
rect -3141 238 -3125 272
rect -3067 238 -3051 272
rect -2883 238 -2867 272
rect -2809 238 -2793 272
rect -2625 238 -2609 272
rect -2551 238 -2535 272
rect -2367 238 -2351 272
rect -2293 238 -2277 272
rect -2109 238 -2093 272
rect -2035 238 -2019 272
rect -1851 238 -1835 272
rect -1777 238 -1761 272
rect -1593 238 -1577 272
rect -1519 238 -1503 272
rect -1335 238 -1319 272
rect -1261 238 -1245 272
rect -1077 238 -1061 272
rect -1003 238 -987 272
rect -819 238 -803 272
rect -745 238 -729 272
rect -561 238 -545 272
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect 545 238 561 272
rect 729 238 745 272
rect 803 238 819 272
rect 987 238 1003 272
rect 1061 238 1077 272
rect 1245 238 1261 272
rect 1319 238 1335 272
rect 1503 238 1519 272
rect 1577 238 1593 272
rect 1761 238 1777 272
rect 1835 238 1851 272
rect 2019 238 2035 272
rect 2093 238 2109 272
rect 2277 238 2293 272
rect 2351 238 2367 272
rect 2535 238 2551 272
rect 2609 238 2625 272
rect 2793 238 2809 272
rect 2867 238 2883 272
rect 3051 238 3067 272
rect 3125 238 3141 272
rect 3309 238 3325 272
rect -3371 188 -3337 204
rect -3371 -204 -3337 -188
rect -3113 188 -3079 204
rect -3113 -204 -3079 -188
rect -2855 188 -2821 204
rect -2855 -204 -2821 -188
rect -2597 188 -2563 204
rect -2597 -204 -2563 -188
rect -2339 188 -2305 204
rect -2339 -204 -2305 -188
rect -2081 188 -2047 204
rect -2081 -204 -2047 -188
rect -1823 188 -1789 204
rect -1823 -204 -1789 -188
rect -1565 188 -1531 204
rect -1565 -204 -1531 -188
rect -1307 188 -1273 204
rect -1307 -204 -1273 -188
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect 1273 188 1307 204
rect 1273 -204 1307 -188
rect 1531 188 1565 204
rect 1531 -204 1565 -188
rect 1789 188 1823 204
rect 1789 -204 1823 -188
rect 2047 188 2081 204
rect 2047 -204 2081 -188
rect 2305 188 2339 204
rect 2305 -204 2339 -188
rect 2563 188 2597 204
rect 2563 -204 2597 -188
rect 2821 188 2855 204
rect 2821 -204 2855 -188
rect 3079 188 3113 204
rect 3079 -204 3113 -188
rect 3337 188 3371 204
rect 3337 -204 3371 -188
rect -3325 -272 -3309 -238
rect -3141 -272 -3125 -238
rect -3067 -272 -3051 -238
rect -2883 -272 -2867 -238
rect -2809 -272 -2793 -238
rect -2625 -272 -2609 -238
rect -2551 -272 -2535 -238
rect -2367 -272 -2351 -238
rect -2293 -272 -2277 -238
rect -2109 -272 -2093 -238
rect -2035 -272 -2019 -238
rect -1851 -272 -1835 -238
rect -1777 -272 -1761 -238
rect -1593 -272 -1577 -238
rect -1519 -272 -1503 -238
rect -1335 -272 -1319 -238
rect -1261 -272 -1245 -238
rect -1077 -272 -1061 -238
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect 1061 -272 1077 -238
rect 1245 -272 1261 -238
rect 1319 -272 1335 -238
rect 1503 -272 1519 -238
rect 1577 -272 1593 -238
rect 1761 -272 1777 -238
rect 1835 -272 1851 -238
rect 2019 -272 2035 -238
rect 2093 -272 2109 -238
rect 2277 -272 2293 -238
rect 2351 -272 2367 -238
rect 2535 -272 2551 -238
rect 2609 -272 2625 -238
rect 2793 -272 2809 -238
rect 2867 -272 2883 -238
rect 3051 -272 3067 -238
rect 3125 -272 3141 -238
rect 3309 -272 3325 -238
rect -3485 -340 -3451 -278
rect 3451 -340 3485 -278
rect -3485 -374 -3389 -340
rect 3389 -374 3485 -340
<< viali >>
rect -3309 238 -3141 272
rect -3051 238 -2883 272
rect -2793 238 -2625 272
rect -2535 238 -2367 272
rect -2277 238 -2109 272
rect -2019 238 -1851 272
rect -1761 238 -1593 272
rect -1503 238 -1335 272
rect -1245 238 -1077 272
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect 1077 238 1245 272
rect 1335 238 1503 272
rect 1593 238 1761 272
rect 1851 238 2019 272
rect 2109 238 2277 272
rect 2367 238 2535 272
rect 2625 238 2793 272
rect 2883 238 3051 272
rect 3141 238 3309 272
rect -3371 -188 -3337 188
rect -3113 -188 -3079 188
rect -2855 -188 -2821 188
rect -2597 -188 -2563 188
rect -2339 -188 -2305 188
rect -2081 -188 -2047 188
rect -1823 -188 -1789 188
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect 1789 -188 1823 188
rect 2047 -188 2081 188
rect 2305 -188 2339 188
rect 2563 -188 2597 188
rect 2821 -188 2855 188
rect 3079 -188 3113 188
rect 3337 -188 3371 188
rect -3309 -272 -3141 -238
rect -3051 -272 -2883 -238
rect -2793 -272 -2625 -238
rect -2535 -272 -2367 -238
rect -2277 -272 -2109 -238
rect -2019 -272 -1851 -238
rect -1761 -272 -1593 -238
rect -1503 -272 -1335 -238
rect -1245 -272 -1077 -238
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
rect 1077 -272 1245 -238
rect 1335 -272 1503 -238
rect 1593 -272 1761 -238
rect 1851 -272 2019 -238
rect 2109 -272 2277 -238
rect 2367 -272 2535 -238
rect 2625 -272 2793 -238
rect 2883 -272 3051 -238
rect 3141 -272 3309 -238
<< metal1 >>
rect -3321 272 -3129 278
rect -3321 238 -3309 272
rect -3141 238 -3129 272
rect -3321 232 -3129 238
rect -3063 272 -2871 278
rect -3063 238 -3051 272
rect -2883 238 -2871 272
rect -3063 232 -2871 238
rect -2805 272 -2613 278
rect -2805 238 -2793 272
rect -2625 238 -2613 272
rect -2805 232 -2613 238
rect -2547 272 -2355 278
rect -2547 238 -2535 272
rect -2367 238 -2355 272
rect -2547 232 -2355 238
rect -2289 272 -2097 278
rect -2289 238 -2277 272
rect -2109 238 -2097 272
rect -2289 232 -2097 238
rect -2031 272 -1839 278
rect -2031 238 -2019 272
rect -1851 238 -1839 272
rect -2031 232 -1839 238
rect -1773 272 -1581 278
rect -1773 238 -1761 272
rect -1593 238 -1581 272
rect -1773 232 -1581 238
rect -1515 272 -1323 278
rect -1515 238 -1503 272
rect -1335 238 -1323 272
rect -1515 232 -1323 238
rect -1257 272 -1065 278
rect -1257 238 -1245 272
rect -1077 238 -1065 272
rect -1257 232 -1065 238
rect -999 272 -807 278
rect -999 238 -987 272
rect -819 238 -807 272
rect -999 232 -807 238
rect -741 272 -549 278
rect -741 238 -729 272
rect -561 238 -549 272
rect -741 232 -549 238
rect -483 272 -291 278
rect -483 238 -471 272
rect -303 238 -291 272
rect -483 232 -291 238
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect 291 272 483 278
rect 291 238 303 272
rect 471 238 483 272
rect 291 232 483 238
rect 549 272 741 278
rect 549 238 561 272
rect 729 238 741 272
rect 549 232 741 238
rect 807 272 999 278
rect 807 238 819 272
rect 987 238 999 272
rect 807 232 999 238
rect 1065 272 1257 278
rect 1065 238 1077 272
rect 1245 238 1257 272
rect 1065 232 1257 238
rect 1323 272 1515 278
rect 1323 238 1335 272
rect 1503 238 1515 272
rect 1323 232 1515 238
rect 1581 272 1773 278
rect 1581 238 1593 272
rect 1761 238 1773 272
rect 1581 232 1773 238
rect 1839 272 2031 278
rect 1839 238 1851 272
rect 2019 238 2031 272
rect 1839 232 2031 238
rect 2097 272 2289 278
rect 2097 238 2109 272
rect 2277 238 2289 272
rect 2097 232 2289 238
rect 2355 272 2547 278
rect 2355 238 2367 272
rect 2535 238 2547 272
rect 2355 232 2547 238
rect 2613 272 2805 278
rect 2613 238 2625 272
rect 2793 238 2805 272
rect 2613 232 2805 238
rect 2871 272 3063 278
rect 2871 238 2883 272
rect 3051 238 3063 272
rect 2871 232 3063 238
rect 3129 272 3321 278
rect 3129 238 3141 272
rect 3309 238 3321 272
rect 3129 232 3321 238
rect -3377 188 -3331 200
rect -3377 -188 -3371 188
rect -3337 -188 -3331 188
rect -3377 -200 -3331 -188
rect -3119 188 -3073 200
rect -3119 -188 -3113 188
rect -3079 -188 -3073 188
rect -3119 -200 -3073 -188
rect -2861 188 -2815 200
rect -2861 -188 -2855 188
rect -2821 -188 -2815 188
rect -2861 -200 -2815 -188
rect -2603 188 -2557 200
rect -2603 -188 -2597 188
rect -2563 -188 -2557 188
rect -2603 -200 -2557 -188
rect -2345 188 -2299 200
rect -2345 -188 -2339 188
rect -2305 -188 -2299 188
rect -2345 -200 -2299 -188
rect -2087 188 -2041 200
rect -2087 -188 -2081 188
rect -2047 -188 -2041 188
rect -2087 -200 -2041 -188
rect -1829 188 -1783 200
rect -1829 -188 -1823 188
rect -1789 -188 -1783 188
rect -1829 -200 -1783 -188
rect -1571 188 -1525 200
rect -1571 -188 -1565 188
rect -1531 -188 -1525 188
rect -1571 -200 -1525 -188
rect -1313 188 -1267 200
rect -1313 -188 -1307 188
rect -1273 -188 -1267 188
rect -1313 -200 -1267 -188
rect -1055 188 -1009 200
rect -1055 -188 -1049 188
rect -1015 -188 -1009 188
rect -1055 -200 -1009 -188
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect 1009 188 1055 200
rect 1009 -188 1015 188
rect 1049 -188 1055 188
rect 1009 -200 1055 -188
rect 1267 188 1313 200
rect 1267 -188 1273 188
rect 1307 -188 1313 188
rect 1267 -200 1313 -188
rect 1525 188 1571 200
rect 1525 -188 1531 188
rect 1565 -188 1571 188
rect 1525 -200 1571 -188
rect 1783 188 1829 200
rect 1783 -188 1789 188
rect 1823 -188 1829 188
rect 1783 -200 1829 -188
rect 2041 188 2087 200
rect 2041 -188 2047 188
rect 2081 -188 2087 188
rect 2041 -200 2087 -188
rect 2299 188 2345 200
rect 2299 -188 2305 188
rect 2339 -188 2345 188
rect 2299 -200 2345 -188
rect 2557 188 2603 200
rect 2557 -188 2563 188
rect 2597 -188 2603 188
rect 2557 -200 2603 -188
rect 2815 188 2861 200
rect 2815 -188 2821 188
rect 2855 -188 2861 188
rect 2815 -200 2861 -188
rect 3073 188 3119 200
rect 3073 -188 3079 188
rect 3113 -188 3119 188
rect 3073 -200 3119 -188
rect 3331 188 3377 200
rect 3331 -188 3337 188
rect 3371 -188 3377 188
rect 3331 -200 3377 -188
rect -3321 -238 -3129 -232
rect -3321 -272 -3309 -238
rect -3141 -272 -3129 -238
rect -3321 -278 -3129 -272
rect -3063 -238 -2871 -232
rect -3063 -272 -3051 -238
rect -2883 -272 -2871 -238
rect -3063 -278 -2871 -272
rect -2805 -238 -2613 -232
rect -2805 -272 -2793 -238
rect -2625 -272 -2613 -238
rect -2805 -278 -2613 -272
rect -2547 -238 -2355 -232
rect -2547 -272 -2535 -238
rect -2367 -272 -2355 -238
rect -2547 -278 -2355 -272
rect -2289 -238 -2097 -232
rect -2289 -272 -2277 -238
rect -2109 -272 -2097 -238
rect -2289 -278 -2097 -272
rect -2031 -238 -1839 -232
rect -2031 -272 -2019 -238
rect -1851 -272 -1839 -238
rect -2031 -278 -1839 -272
rect -1773 -238 -1581 -232
rect -1773 -272 -1761 -238
rect -1593 -272 -1581 -238
rect -1773 -278 -1581 -272
rect -1515 -238 -1323 -232
rect -1515 -272 -1503 -238
rect -1335 -272 -1323 -238
rect -1515 -278 -1323 -272
rect -1257 -238 -1065 -232
rect -1257 -272 -1245 -238
rect -1077 -272 -1065 -238
rect -1257 -278 -1065 -272
rect -999 -238 -807 -232
rect -999 -272 -987 -238
rect -819 -272 -807 -238
rect -999 -278 -807 -272
rect -741 -238 -549 -232
rect -741 -272 -729 -238
rect -561 -272 -549 -238
rect -741 -278 -549 -272
rect -483 -238 -291 -232
rect -483 -272 -471 -238
rect -303 -272 -291 -238
rect -483 -278 -291 -272
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
rect 291 -238 483 -232
rect 291 -272 303 -238
rect 471 -272 483 -238
rect 291 -278 483 -272
rect 549 -238 741 -232
rect 549 -272 561 -238
rect 729 -272 741 -238
rect 549 -278 741 -272
rect 807 -238 999 -232
rect 807 -272 819 -238
rect 987 -272 999 -238
rect 807 -278 999 -272
rect 1065 -238 1257 -232
rect 1065 -272 1077 -238
rect 1245 -272 1257 -238
rect 1065 -278 1257 -272
rect 1323 -238 1515 -232
rect 1323 -272 1335 -238
rect 1503 -272 1515 -238
rect 1323 -278 1515 -272
rect 1581 -238 1773 -232
rect 1581 -272 1593 -238
rect 1761 -272 1773 -238
rect 1581 -278 1773 -272
rect 1839 -238 2031 -232
rect 1839 -272 1851 -238
rect 2019 -272 2031 -238
rect 1839 -278 2031 -272
rect 2097 -238 2289 -232
rect 2097 -272 2109 -238
rect 2277 -272 2289 -238
rect 2097 -278 2289 -272
rect 2355 -238 2547 -232
rect 2355 -272 2367 -238
rect 2535 -272 2547 -238
rect 2355 -278 2547 -272
rect 2613 -238 2805 -232
rect 2613 -272 2625 -238
rect 2793 -272 2805 -238
rect 2613 -278 2805 -272
rect 2871 -238 3063 -232
rect 2871 -272 2883 -238
rect 3051 -272 3063 -238
rect 2871 -278 3063 -272
rect 3129 -238 3321 -232
rect 3129 -272 3141 -238
rect 3309 -272 3321 -238
rect 3129 -278 3321 -272
<< properties >>
string FIXED_BBOX -3468 -357 3468 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
