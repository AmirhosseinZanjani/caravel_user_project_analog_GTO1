magic
tech sky130A
magscale 1 2
timestamp 1698055914
<< nwell >>
rect -16631 -3919 16631 3919
<< pmos >>
rect -16435 -3700 -14435 3700
rect -14377 -3700 -12377 3700
rect -12319 -3700 -10319 3700
rect -10261 -3700 -8261 3700
rect -8203 -3700 -6203 3700
rect -6145 -3700 -4145 3700
rect -4087 -3700 -2087 3700
rect -2029 -3700 -29 3700
rect 29 -3700 2029 3700
rect 2087 -3700 4087 3700
rect 4145 -3700 6145 3700
rect 6203 -3700 8203 3700
rect 8261 -3700 10261 3700
rect 10319 -3700 12319 3700
rect 12377 -3700 14377 3700
rect 14435 -3700 16435 3700
<< pdiff >>
rect -16493 3688 -16435 3700
rect -16493 -3688 -16481 3688
rect -16447 -3688 -16435 3688
rect -16493 -3700 -16435 -3688
rect -14435 3688 -14377 3700
rect -14435 -3688 -14423 3688
rect -14389 -3688 -14377 3688
rect -14435 -3700 -14377 -3688
rect -12377 3688 -12319 3700
rect -12377 -3688 -12365 3688
rect -12331 -3688 -12319 3688
rect -12377 -3700 -12319 -3688
rect -10319 3688 -10261 3700
rect -10319 -3688 -10307 3688
rect -10273 -3688 -10261 3688
rect -10319 -3700 -10261 -3688
rect -8261 3688 -8203 3700
rect -8261 -3688 -8249 3688
rect -8215 -3688 -8203 3688
rect -8261 -3700 -8203 -3688
rect -6203 3688 -6145 3700
rect -6203 -3688 -6191 3688
rect -6157 -3688 -6145 3688
rect -6203 -3700 -6145 -3688
rect -4145 3688 -4087 3700
rect -4145 -3688 -4133 3688
rect -4099 -3688 -4087 3688
rect -4145 -3700 -4087 -3688
rect -2087 3688 -2029 3700
rect -2087 -3688 -2075 3688
rect -2041 -3688 -2029 3688
rect -2087 -3700 -2029 -3688
rect -29 3688 29 3700
rect -29 -3688 -17 3688
rect 17 -3688 29 3688
rect -29 -3700 29 -3688
rect 2029 3688 2087 3700
rect 2029 -3688 2041 3688
rect 2075 -3688 2087 3688
rect 2029 -3700 2087 -3688
rect 4087 3688 4145 3700
rect 4087 -3688 4099 3688
rect 4133 -3688 4145 3688
rect 4087 -3700 4145 -3688
rect 6145 3688 6203 3700
rect 6145 -3688 6157 3688
rect 6191 -3688 6203 3688
rect 6145 -3700 6203 -3688
rect 8203 3688 8261 3700
rect 8203 -3688 8215 3688
rect 8249 -3688 8261 3688
rect 8203 -3700 8261 -3688
rect 10261 3688 10319 3700
rect 10261 -3688 10273 3688
rect 10307 -3688 10319 3688
rect 10261 -3700 10319 -3688
rect 12319 3688 12377 3700
rect 12319 -3688 12331 3688
rect 12365 -3688 12377 3688
rect 12319 -3700 12377 -3688
rect 14377 3688 14435 3700
rect 14377 -3688 14389 3688
rect 14423 -3688 14435 3688
rect 14377 -3700 14435 -3688
rect 16435 3688 16493 3700
rect 16435 -3688 16447 3688
rect 16481 -3688 16493 3688
rect 16435 -3700 16493 -3688
<< pdiffc >>
rect -16481 -3688 -16447 3688
rect -14423 -3688 -14389 3688
rect -12365 -3688 -12331 3688
rect -10307 -3688 -10273 3688
rect -8249 -3688 -8215 3688
rect -6191 -3688 -6157 3688
rect -4133 -3688 -4099 3688
rect -2075 -3688 -2041 3688
rect -17 -3688 17 3688
rect 2041 -3688 2075 3688
rect 4099 -3688 4133 3688
rect 6157 -3688 6191 3688
rect 8215 -3688 8249 3688
rect 10273 -3688 10307 3688
rect 12331 -3688 12365 3688
rect 14389 -3688 14423 3688
rect 16447 -3688 16481 3688
<< nsubdiff >>
rect -16595 3849 -16499 3883
rect 16499 3849 16595 3883
rect -16595 3787 -16561 3849
rect 16561 3787 16595 3849
rect -16595 -3849 -16561 -3787
rect 16561 -3849 16595 -3787
rect -16595 -3883 -16499 -3849
rect 16499 -3883 16595 -3849
<< nsubdiffcont >>
rect -16499 3849 16499 3883
rect -16595 -3787 -16561 3787
rect 16561 -3787 16595 3787
rect -16499 -3883 16499 -3849
<< poly >>
rect -16435 3781 -14435 3797
rect -16435 3747 -16419 3781
rect -14451 3747 -14435 3781
rect -16435 3700 -14435 3747
rect -14377 3781 -12377 3797
rect -14377 3747 -14361 3781
rect -12393 3747 -12377 3781
rect -14377 3700 -12377 3747
rect -12319 3781 -10319 3797
rect -12319 3747 -12303 3781
rect -10335 3747 -10319 3781
rect -12319 3700 -10319 3747
rect -10261 3781 -8261 3797
rect -10261 3747 -10245 3781
rect -8277 3747 -8261 3781
rect -10261 3700 -8261 3747
rect -8203 3781 -6203 3797
rect -8203 3747 -8187 3781
rect -6219 3747 -6203 3781
rect -8203 3700 -6203 3747
rect -6145 3781 -4145 3797
rect -6145 3747 -6129 3781
rect -4161 3747 -4145 3781
rect -6145 3700 -4145 3747
rect -4087 3781 -2087 3797
rect -4087 3747 -4071 3781
rect -2103 3747 -2087 3781
rect -4087 3700 -2087 3747
rect -2029 3781 -29 3797
rect -2029 3747 -2013 3781
rect -45 3747 -29 3781
rect -2029 3700 -29 3747
rect 29 3781 2029 3797
rect 29 3747 45 3781
rect 2013 3747 2029 3781
rect 29 3700 2029 3747
rect 2087 3781 4087 3797
rect 2087 3747 2103 3781
rect 4071 3747 4087 3781
rect 2087 3700 4087 3747
rect 4145 3781 6145 3797
rect 4145 3747 4161 3781
rect 6129 3747 6145 3781
rect 4145 3700 6145 3747
rect 6203 3781 8203 3797
rect 6203 3747 6219 3781
rect 8187 3747 8203 3781
rect 6203 3700 8203 3747
rect 8261 3781 10261 3797
rect 8261 3747 8277 3781
rect 10245 3747 10261 3781
rect 8261 3700 10261 3747
rect 10319 3781 12319 3797
rect 10319 3747 10335 3781
rect 12303 3747 12319 3781
rect 10319 3700 12319 3747
rect 12377 3781 14377 3797
rect 12377 3747 12393 3781
rect 14361 3747 14377 3781
rect 12377 3700 14377 3747
rect 14435 3781 16435 3797
rect 14435 3747 14451 3781
rect 16419 3747 16435 3781
rect 14435 3700 16435 3747
rect -16435 -3747 -14435 -3700
rect -16435 -3781 -16419 -3747
rect -14451 -3781 -14435 -3747
rect -16435 -3797 -14435 -3781
rect -14377 -3747 -12377 -3700
rect -14377 -3781 -14361 -3747
rect -12393 -3781 -12377 -3747
rect -14377 -3797 -12377 -3781
rect -12319 -3747 -10319 -3700
rect -12319 -3781 -12303 -3747
rect -10335 -3781 -10319 -3747
rect -12319 -3797 -10319 -3781
rect -10261 -3747 -8261 -3700
rect -10261 -3781 -10245 -3747
rect -8277 -3781 -8261 -3747
rect -10261 -3797 -8261 -3781
rect -8203 -3747 -6203 -3700
rect -8203 -3781 -8187 -3747
rect -6219 -3781 -6203 -3747
rect -8203 -3797 -6203 -3781
rect -6145 -3747 -4145 -3700
rect -6145 -3781 -6129 -3747
rect -4161 -3781 -4145 -3747
rect -6145 -3797 -4145 -3781
rect -4087 -3747 -2087 -3700
rect -4087 -3781 -4071 -3747
rect -2103 -3781 -2087 -3747
rect -4087 -3797 -2087 -3781
rect -2029 -3747 -29 -3700
rect -2029 -3781 -2013 -3747
rect -45 -3781 -29 -3747
rect -2029 -3797 -29 -3781
rect 29 -3747 2029 -3700
rect 29 -3781 45 -3747
rect 2013 -3781 2029 -3747
rect 29 -3797 2029 -3781
rect 2087 -3747 4087 -3700
rect 2087 -3781 2103 -3747
rect 4071 -3781 4087 -3747
rect 2087 -3797 4087 -3781
rect 4145 -3747 6145 -3700
rect 4145 -3781 4161 -3747
rect 6129 -3781 6145 -3747
rect 4145 -3797 6145 -3781
rect 6203 -3747 8203 -3700
rect 6203 -3781 6219 -3747
rect 8187 -3781 8203 -3747
rect 6203 -3797 8203 -3781
rect 8261 -3747 10261 -3700
rect 8261 -3781 8277 -3747
rect 10245 -3781 10261 -3747
rect 8261 -3797 10261 -3781
rect 10319 -3747 12319 -3700
rect 10319 -3781 10335 -3747
rect 12303 -3781 12319 -3747
rect 10319 -3797 12319 -3781
rect 12377 -3747 14377 -3700
rect 12377 -3781 12393 -3747
rect 14361 -3781 14377 -3747
rect 12377 -3797 14377 -3781
rect 14435 -3747 16435 -3700
rect 14435 -3781 14451 -3747
rect 16419 -3781 16435 -3747
rect 14435 -3797 16435 -3781
<< polycont >>
rect -16419 3747 -14451 3781
rect -14361 3747 -12393 3781
rect -12303 3747 -10335 3781
rect -10245 3747 -8277 3781
rect -8187 3747 -6219 3781
rect -6129 3747 -4161 3781
rect -4071 3747 -2103 3781
rect -2013 3747 -45 3781
rect 45 3747 2013 3781
rect 2103 3747 4071 3781
rect 4161 3747 6129 3781
rect 6219 3747 8187 3781
rect 8277 3747 10245 3781
rect 10335 3747 12303 3781
rect 12393 3747 14361 3781
rect 14451 3747 16419 3781
rect -16419 -3781 -14451 -3747
rect -14361 -3781 -12393 -3747
rect -12303 -3781 -10335 -3747
rect -10245 -3781 -8277 -3747
rect -8187 -3781 -6219 -3747
rect -6129 -3781 -4161 -3747
rect -4071 -3781 -2103 -3747
rect -2013 -3781 -45 -3747
rect 45 -3781 2013 -3747
rect 2103 -3781 4071 -3747
rect 4161 -3781 6129 -3747
rect 6219 -3781 8187 -3747
rect 8277 -3781 10245 -3747
rect 10335 -3781 12303 -3747
rect 12393 -3781 14361 -3747
rect 14451 -3781 16419 -3747
<< locali >>
rect -16595 3849 -16499 3883
rect 16499 3849 16595 3883
rect -16595 3787 -16561 3849
rect 16561 3787 16595 3849
rect -16435 3747 -16419 3781
rect -14451 3747 -14435 3781
rect -14377 3747 -14361 3781
rect -12393 3747 -12377 3781
rect -12319 3747 -12303 3781
rect -10335 3747 -10319 3781
rect -10261 3747 -10245 3781
rect -8277 3747 -8261 3781
rect -8203 3747 -8187 3781
rect -6219 3747 -6203 3781
rect -6145 3747 -6129 3781
rect -4161 3747 -4145 3781
rect -4087 3747 -4071 3781
rect -2103 3747 -2087 3781
rect -2029 3747 -2013 3781
rect -45 3747 -29 3781
rect 29 3747 45 3781
rect 2013 3747 2029 3781
rect 2087 3747 2103 3781
rect 4071 3747 4087 3781
rect 4145 3747 4161 3781
rect 6129 3747 6145 3781
rect 6203 3747 6219 3781
rect 8187 3747 8203 3781
rect 8261 3747 8277 3781
rect 10245 3747 10261 3781
rect 10319 3747 10335 3781
rect 12303 3747 12319 3781
rect 12377 3747 12393 3781
rect 14361 3747 14377 3781
rect 14435 3747 14451 3781
rect 16419 3747 16435 3781
rect -16481 3688 -16447 3704
rect -16481 -3704 -16447 -3688
rect -14423 3688 -14389 3704
rect -14423 -3704 -14389 -3688
rect -12365 3688 -12331 3704
rect -12365 -3704 -12331 -3688
rect -10307 3688 -10273 3704
rect -10307 -3704 -10273 -3688
rect -8249 3688 -8215 3704
rect -8249 -3704 -8215 -3688
rect -6191 3688 -6157 3704
rect -6191 -3704 -6157 -3688
rect -4133 3688 -4099 3704
rect -4133 -3704 -4099 -3688
rect -2075 3688 -2041 3704
rect -2075 -3704 -2041 -3688
rect -17 3688 17 3704
rect -17 -3704 17 -3688
rect 2041 3688 2075 3704
rect 2041 -3704 2075 -3688
rect 4099 3688 4133 3704
rect 4099 -3704 4133 -3688
rect 6157 3688 6191 3704
rect 6157 -3704 6191 -3688
rect 8215 3688 8249 3704
rect 8215 -3704 8249 -3688
rect 10273 3688 10307 3704
rect 10273 -3704 10307 -3688
rect 12331 3688 12365 3704
rect 12331 -3704 12365 -3688
rect 14389 3688 14423 3704
rect 14389 -3704 14423 -3688
rect 16447 3688 16481 3704
rect 16447 -3704 16481 -3688
rect -16435 -3781 -16419 -3747
rect -14451 -3781 -14435 -3747
rect -14377 -3781 -14361 -3747
rect -12393 -3781 -12377 -3747
rect -12319 -3781 -12303 -3747
rect -10335 -3781 -10319 -3747
rect -10261 -3781 -10245 -3747
rect -8277 -3781 -8261 -3747
rect -8203 -3781 -8187 -3747
rect -6219 -3781 -6203 -3747
rect -6145 -3781 -6129 -3747
rect -4161 -3781 -4145 -3747
rect -4087 -3781 -4071 -3747
rect -2103 -3781 -2087 -3747
rect -2029 -3781 -2013 -3747
rect -45 -3781 -29 -3747
rect 29 -3781 45 -3747
rect 2013 -3781 2029 -3747
rect 2087 -3781 2103 -3747
rect 4071 -3781 4087 -3747
rect 4145 -3781 4161 -3747
rect 6129 -3781 6145 -3747
rect 6203 -3781 6219 -3747
rect 8187 -3781 8203 -3747
rect 8261 -3781 8277 -3747
rect 10245 -3781 10261 -3747
rect 10319 -3781 10335 -3747
rect 12303 -3781 12319 -3747
rect 12377 -3781 12393 -3747
rect 14361 -3781 14377 -3747
rect 14435 -3781 14451 -3747
rect 16419 -3781 16435 -3747
rect -16595 -3849 -16561 -3787
rect 16561 -3849 16595 -3787
rect -16595 -3883 -16499 -3849
rect 16499 -3883 16595 -3849
<< viali >>
rect -16419 3747 -14451 3781
rect -14361 3747 -12393 3781
rect -12303 3747 -10335 3781
rect -10245 3747 -8277 3781
rect -8187 3747 -6219 3781
rect -6129 3747 -4161 3781
rect -4071 3747 -2103 3781
rect -2013 3747 -45 3781
rect 45 3747 2013 3781
rect 2103 3747 4071 3781
rect 4161 3747 6129 3781
rect 6219 3747 8187 3781
rect 8277 3747 10245 3781
rect 10335 3747 12303 3781
rect 12393 3747 14361 3781
rect 14451 3747 16419 3781
rect -16481 -3688 -16447 3688
rect -14423 -3688 -14389 3688
rect -12365 -3688 -12331 3688
rect -10307 -3688 -10273 3688
rect -8249 -3688 -8215 3688
rect -6191 -3688 -6157 3688
rect -4133 -3688 -4099 3688
rect -2075 -3688 -2041 3688
rect -17 -3688 17 3688
rect 2041 -3688 2075 3688
rect 4099 -3688 4133 3688
rect 6157 -3688 6191 3688
rect 8215 -3688 8249 3688
rect 10273 -3688 10307 3688
rect 12331 -3688 12365 3688
rect 14389 -3688 14423 3688
rect 16447 -3688 16481 3688
rect -16419 -3781 -14451 -3747
rect -14361 -3781 -12393 -3747
rect -12303 -3781 -10335 -3747
rect -10245 -3781 -8277 -3747
rect -8187 -3781 -6219 -3747
rect -6129 -3781 -4161 -3747
rect -4071 -3781 -2103 -3747
rect -2013 -3781 -45 -3747
rect 45 -3781 2013 -3747
rect 2103 -3781 4071 -3747
rect 4161 -3781 6129 -3747
rect 6219 -3781 8187 -3747
rect 8277 -3781 10245 -3747
rect 10335 -3781 12303 -3747
rect 12393 -3781 14361 -3747
rect 14451 -3781 16419 -3747
<< metal1 >>
rect -16431 3781 -14439 3787
rect -16431 3747 -16419 3781
rect -14451 3747 -14439 3781
rect -16431 3741 -14439 3747
rect -14373 3781 -12381 3787
rect -14373 3747 -14361 3781
rect -12393 3747 -12381 3781
rect -14373 3741 -12381 3747
rect -12315 3781 -10323 3787
rect -12315 3747 -12303 3781
rect -10335 3747 -10323 3781
rect -12315 3741 -10323 3747
rect -10257 3781 -8265 3787
rect -10257 3747 -10245 3781
rect -8277 3747 -8265 3781
rect -10257 3741 -8265 3747
rect -8199 3781 -6207 3787
rect -8199 3747 -8187 3781
rect -6219 3747 -6207 3781
rect -8199 3741 -6207 3747
rect -6141 3781 -4149 3787
rect -6141 3747 -6129 3781
rect -4161 3747 -4149 3781
rect -6141 3741 -4149 3747
rect -4083 3781 -2091 3787
rect -4083 3747 -4071 3781
rect -2103 3747 -2091 3781
rect -4083 3741 -2091 3747
rect -2025 3781 -33 3787
rect -2025 3747 -2013 3781
rect -45 3747 -33 3781
rect -2025 3741 -33 3747
rect 33 3781 2025 3787
rect 33 3747 45 3781
rect 2013 3747 2025 3781
rect 33 3741 2025 3747
rect 2091 3781 4083 3787
rect 2091 3747 2103 3781
rect 4071 3747 4083 3781
rect 2091 3741 4083 3747
rect 4149 3781 6141 3787
rect 4149 3747 4161 3781
rect 6129 3747 6141 3781
rect 4149 3741 6141 3747
rect 6207 3781 8199 3787
rect 6207 3747 6219 3781
rect 8187 3747 8199 3781
rect 6207 3741 8199 3747
rect 8265 3781 10257 3787
rect 8265 3747 8277 3781
rect 10245 3747 10257 3781
rect 8265 3741 10257 3747
rect 10323 3781 12315 3787
rect 10323 3747 10335 3781
rect 12303 3747 12315 3781
rect 10323 3741 12315 3747
rect 12381 3781 14373 3787
rect 12381 3747 12393 3781
rect 14361 3747 14373 3781
rect 12381 3741 14373 3747
rect 14439 3781 16431 3787
rect 14439 3747 14451 3781
rect 16419 3747 16431 3781
rect 14439 3741 16431 3747
rect -16487 3688 -16441 3700
rect -16487 -3688 -16481 3688
rect -16447 -3688 -16441 3688
rect -16487 -3700 -16441 -3688
rect -14429 3688 -14383 3700
rect -14429 -3688 -14423 3688
rect -14389 -3688 -14383 3688
rect -14429 -3700 -14383 -3688
rect -12371 3688 -12325 3700
rect -12371 -3688 -12365 3688
rect -12331 -3688 -12325 3688
rect -12371 -3700 -12325 -3688
rect -10313 3688 -10267 3700
rect -10313 -3688 -10307 3688
rect -10273 -3688 -10267 3688
rect -10313 -3700 -10267 -3688
rect -8255 3688 -8209 3700
rect -8255 -3688 -8249 3688
rect -8215 -3688 -8209 3688
rect -8255 -3700 -8209 -3688
rect -6197 3688 -6151 3700
rect -6197 -3688 -6191 3688
rect -6157 -3688 -6151 3688
rect -6197 -3700 -6151 -3688
rect -4139 3688 -4093 3700
rect -4139 -3688 -4133 3688
rect -4099 -3688 -4093 3688
rect -4139 -3700 -4093 -3688
rect -2081 3688 -2035 3700
rect -2081 -3688 -2075 3688
rect -2041 -3688 -2035 3688
rect -2081 -3700 -2035 -3688
rect -23 3688 23 3700
rect -23 -3688 -17 3688
rect 17 -3688 23 3688
rect -23 -3700 23 -3688
rect 2035 3688 2081 3700
rect 2035 -3688 2041 3688
rect 2075 -3688 2081 3688
rect 2035 -3700 2081 -3688
rect 4093 3688 4139 3700
rect 4093 -3688 4099 3688
rect 4133 -3688 4139 3688
rect 4093 -3700 4139 -3688
rect 6151 3688 6197 3700
rect 6151 -3688 6157 3688
rect 6191 -3688 6197 3688
rect 6151 -3700 6197 -3688
rect 8209 3688 8255 3700
rect 8209 -3688 8215 3688
rect 8249 -3688 8255 3688
rect 8209 -3700 8255 -3688
rect 10267 3688 10313 3700
rect 10267 -3688 10273 3688
rect 10307 -3688 10313 3688
rect 10267 -3700 10313 -3688
rect 12325 3688 12371 3700
rect 12325 -3688 12331 3688
rect 12365 -3688 12371 3688
rect 12325 -3700 12371 -3688
rect 14383 3688 14429 3700
rect 14383 -3688 14389 3688
rect 14423 -3688 14429 3688
rect 14383 -3700 14429 -3688
rect 16441 3688 16487 3700
rect 16441 -3688 16447 3688
rect 16481 -3688 16487 3688
rect 16441 -3700 16487 -3688
rect -16431 -3747 -14439 -3741
rect -16431 -3781 -16419 -3747
rect -14451 -3781 -14439 -3747
rect -16431 -3787 -14439 -3781
rect -14373 -3747 -12381 -3741
rect -14373 -3781 -14361 -3747
rect -12393 -3781 -12381 -3747
rect -14373 -3787 -12381 -3781
rect -12315 -3747 -10323 -3741
rect -12315 -3781 -12303 -3747
rect -10335 -3781 -10323 -3747
rect -12315 -3787 -10323 -3781
rect -10257 -3747 -8265 -3741
rect -10257 -3781 -10245 -3747
rect -8277 -3781 -8265 -3747
rect -10257 -3787 -8265 -3781
rect -8199 -3747 -6207 -3741
rect -8199 -3781 -8187 -3747
rect -6219 -3781 -6207 -3747
rect -8199 -3787 -6207 -3781
rect -6141 -3747 -4149 -3741
rect -6141 -3781 -6129 -3747
rect -4161 -3781 -4149 -3747
rect -6141 -3787 -4149 -3781
rect -4083 -3747 -2091 -3741
rect -4083 -3781 -4071 -3747
rect -2103 -3781 -2091 -3747
rect -4083 -3787 -2091 -3781
rect -2025 -3747 -33 -3741
rect -2025 -3781 -2013 -3747
rect -45 -3781 -33 -3747
rect -2025 -3787 -33 -3781
rect 33 -3747 2025 -3741
rect 33 -3781 45 -3747
rect 2013 -3781 2025 -3747
rect 33 -3787 2025 -3781
rect 2091 -3747 4083 -3741
rect 2091 -3781 2103 -3747
rect 4071 -3781 4083 -3747
rect 2091 -3787 4083 -3781
rect 4149 -3747 6141 -3741
rect 4149 -3781 4161 -3747
rect 6129 -3781 6141 -3747
rect 4149 -3787 6141 -3781
rect 6207 -3747 8199 -3741
rect 6207 -3781 6219 -3747
rect 8187 -3781 8199 -3747
rect 6207 -3787 8199 -3781
rect 8265 -3747 10257 -3741
rect 8265 -3781 8277 -3747
rect 10245 -3781 10257 -3747
rect 8265 -3787 10257 -3781
rect 10323 -3747 12315 -3741
rect 10323 -3781 10335 -3747
rect 12303 -3781 12315 -3747
rect 10323 -3787 12315 -3781
rect 12381 -3747 14373 -3741
rect 12381 -3781 12393 -3747
rect 14361 -3781 14373 -3747
rect 12381 -3787 14373 -3781
rect 14439 -3747 16431 -3741
rect 14439 -3781 14451 -3747
rect 16419 -3781 16431 -3747
rect 14439 -3787 16431 -3781
<< properties >>
string FIXED_BBOX -16578 -3866 16578 3866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 37 l 10 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
