magic
tech sky130A
magscale 1 2
timestamp 1693401401
<< error_p >>
rect -941 114 -883 120
rect -749 114 -691 120
rect -557 114 -499 120
rect -365 114 -307 120
rect -173 114 -115 120
rect 19 114 77 120
rect 211 114 269 120
rect 403 114 461 120
rect 595 114 653 120
rect 787 114 845 120
rect 979 114 1037 120
rect -941 80 -929 114
rect -749 80 -737 114
rect -557 80 -545 114
rect -365 80 -353 114
rect -173 80 -161 114
rect 19 80 31 114
rect 211 80 223 114
rect 403 80 415 114
rect 595 80 607 114
rect 787 80 799 114
rect 979 80 991 114
rect -941 74 -883 80
rect -749 74 -691 80
rect -557 74 -499 80
rect -365 74 -307 80
rect -173 74 -115 80
rect 19 74 77 80
rect 211 74 269 80
rect 403 74 461 80
rect 595 74 653 80
rect 787 74 845 80
rect 979 74 1037 80
rect -1037 -80 -979 -74
rect -845 -80 -787 -74
rect -653 -80 -595 -74
rect -461 -80 -403 -74
rect -269 -80 -211 -74
rect -77 -80 -19 -74
rect 115 -80 173 -74
rect 307 -80 365 -74
rect 499 -80 557 -74
rect 691 -80 749 -74
rect 883 -80 941 -74
rect -1037 -114 -1025 -80
rect -845 -114 -833 -80
rect -653 -114 -641 -80
rect -461 -114 -449 -80
rect -269 -114 -257 -80
rect -77 -114 -65 -80
rect 115 -114 127 -80
rect 307 -114 319 -80
rect 499 -114 511 -80
rect 691 -114 703 -80
rect 883 -114 895 -80
rect -1037 -120 -979 -114
rect -845 -120 -787 -114
rect -653 -120 -595 -114
rect -461 -120 -403 -114
rect -269 -120 -211 -114
rect -77 -120 -19 -114
rect 115 -120 173 -114
rect 307 -120 365 -114
rect 499 -120 557 -114
rect 691 -120 749 -114
rect 883 -120 941 -114
<< pwell >>
rect -1223 -252 1223 252
<< nmos >>
rect -1023 -42 -993 42
rect -927 -42 -897 42
rect -831 -42 -801 42
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
rect 801 -42 831 42
rect 897 -42 927 42
rect 993 -42 1023 42
<< ndiff >>
rect -1085 30 -1023 42
rect -1085 -30 -1073 30
rect -1039 -30 -1023 30
rect -1085 -42 -1023 -30
rect -993 30 -927 42
rect -993 -30 -977 30
rect -943 -30 -927 30
rect -993 -42 -927 -30
rect -897 30 -831 42
rect -897 -30 -881 30
rect -847 -30 -831 30
rect -897 -42 -831 -30
rect -801 30 -735 42
rect -801 -30 -785 30
rect -751 -30 -735 30
rect -801 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 801 42
rect 735 -30 751 30
rect 785 -30 801 30
rect 735 -42 801 -30
rect 831 30 897 42
rect 831 -30 847 30
rect 881 -30 897 30
rect 831 -42 897 -30
rect 927 30 993 42
rect 927 -30 943 30
rect 977 -30 993 30
rect 927 -42 993 -30
rect 1023 30 1085 42
rect 1023 -30 1039 30
rect 1073 -30 1085 30
rect 1023 -42 1085 -30
<< ndiffc >>
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
<< psubdiff >>
rect -1187 182 -1091 216
rect 1091 182 1187 216
rect -1187 120 -1153 182
rect 1153 120 1187 182
rect -1187 -182 -1153 -120
rect 1153 -182 1187 -120
rect -1187 -216 -1091 -182
rect 1091 -216 1187 -182
<< psubdiffcont >>
rect -1091 182 1091 216
rect -1187 -120 -1153 120
rect 1153 -120 1187 120
rect -1091 -216 1091 -182
<< poly >>
rect -945 114 -879 130
rect -945 80 -929 114
rect -895 80 -879 114
rect -1023 42 -993 68
rect -945 64 -879 80
rect -753 114 -687 130
rect -753 80 -737 114
rect -703 80 -687 114
rect -927 42 -897 64
rect -831 42 -801 68
rect -753 64 -687 80
rect -561 114 -495 130
rect -561 80 -545 114
rect -511 80 -495 114
rect -735 42 -705 64
rect -639 42 -609 68
rect -561 64 -495 80
rect -369 114 -303 130
rect -369 80 -353 114
rect -319 80 -303 114
rect -543 42 -513 64
rect -447 42 -417 68
rect -369 64 -303 80
rect -177 114 -111 130
rect -177 80 -161 114
rect -127 80 -111 114
rect -351 42 -321 64
rect -255 42 -225 68
rect -177 64 -111 80
rect 15 114 81 130
rect 15 80 31 114
rect 65 80 81 114
rect -159 42 -129 64
rect -63 42 -33 68
rect 15 64 81 80
rect 207 114 273 130
rect 207 80 223 114
rect 257 80 273 114
rect 33 42 63 64
rect 129 42 159 68
rect 207 64 273 80
rect 399 114 465 130
rect 399 80 415 114
rect 449 80 465 114
rect 225 42 255 64
rect 321 42 351 68
rect 399 64 465 80
rect 591 114 657 130
rect 591 80 607 114
rect 641 80 657 114
rect 417 42 447 64
rect 513 42 543 68
rect 591 64 657 80
rect 783 114 849 130
rect 783 80 799 114
rect 833 80 849 114
rect 609 42 639 64
rect 705 42 735 68
rect 783 64 849 80
rect 975 114 1041 130
rect 975 80 991 114
rect 1025 80 1041 114
rect 801 42 831 64
rect 897 42 927 68
rect 975 64 1041 80
rect 993 42 1023 64
rect -1023 -64 -993 -42
rect -1041 -80 -975 -64
rect -927 -68 -897 -42
rect -831 -64 -801 -42
rect -1041 -114 -1025 -80
rect -991 -114 -975 -80
rect -1041 -130 -975 -114
rect -849 -80 -783 -64
rect -735 -68 -705 -42
rect -639 -64 -609 -42
rect -849 -114 -833 -80
rect -799 -114 -783 -80
rect -849 -130 -783 -114
rect -657 -80 -591 -64
rect -543 -68 -513 -42
rect -447 -64 -417 -42
rect -657 -114 -641 -80
rect -607 -114 -591 -80
rect -657 -130 -591 -114
rect -465 -80 -399 -64
rect -351 -68 -321 -42
rect -255 -64 -225 -42
rect -465 -114 -449 -80
rect -415 -114 -399 -80
rect -465 -130 -399 -114
rect -273 -80 -207 -64
rect -159 -68 -129 -42
rect -63 -64 -33 -42
rect -273 -114 -257 -80
rect -223 -114 -207 -80
rect -273 -130 -207 -114
rect -81 -80 -15 -64
rect 33 -68 63 -42
rect 129 -64 159 -42
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect -81 -130 -15 -114
rect 111 -80 177 -64
rect 225 -68 255 -42
rect 321 -64 351 -42
rect 111 -114 127 -80
rect 161 -114 177 -80
rect 111 -130 177 -114
rect 303 -80 369 -64
rect 417 -68 447 -42
rect 513 -64 543 -42
rect 303 -114 319 -80
rect 353 -114 369 -80
rect 303 -130 369 -114
rect 495 -80 561 -64
rect 609 -68 639 -42
rect 705 -64 735 -42
rect 495 -114 511 -80
rect 545 -114 561 -80
rect 495 -130 561 -114
rect 687 -80 753 -64
rect 801 -68 831 -42
rect 897 -64 927 -42
rect 687 -114 703 -80
rect 737 -114 753 -80
rect 687 -130 753 -114
rect 879 -80 945 -64
rect 993 -68 1023 -42
rect 879 -114 895 -80
rect 929 -114 945 -80
rect 879 -130 945 -114
<< polycont >>
rect -929 80 -895 114
rect -737 80 -703 114
rect -545 80 -511 114
rect -353 80 -319 114
rect -161 80 -127 114
rect 31 80 65 114
rect 223 80 257 114
rect 415 80 449 114
rect 607 80 641 114
rect 799 80 833 114
rect 991 80 1025 114
rect -1025 -114 -991 -80
rect -833 -114 -799 -80
rect -641 -114 -607 -80
rect -449 -114 -415 -80
rect -257 -114 -223 -80
rect -65 -114 -31 -80
rect 127 -114 161 -80
rect 319 -114 353 -80
rect 511 -114 545 -80
rect 703 -114 737 -80
rect 895 -114 929 -80
<< locali >>
rect -1187 182 -1091 216
rect 1091 182 1187 216
rect -1187 120 -1153 182
rect 1153 120 1187 182
rect -945 80 -929 114
rect -895 80 -879 114
rect -753 80 -737 114
rect -703 80 -687 114
rect -561 80 -545 114
rect -511 80 -495 114
rect -369 80 -353 114
rect -319 80 -303 114
rect -177 80 -161 114
rect -127 80 -111 114
rect 15 80 31 114
rect 65 80 81 114
rect 207 80 223 114
rect 257 80 273 114
rect 399 80 415 114
rect 449 80 465 114
rect 591 80 607 114
rect 641 80 657 114
rect 783 80 799 114
rect 833 80 849 114
rect 975 80 991 114
rect 1025 80 1041 114
rect -1073 30 -1039 46
rect -1073 -46 -1039 -30
rect -977 30 -943 46
rect -977 -46 -943 -30
rect -881 30 -847 46
rect -881 -46 -847 -30
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect 847 30 881 46
rect 847 -46 881 -30
rect 943 30 977 46
rect 943 -46 977 -30
rect 1039 30 1073 46
rect 1039 -46 1073 -30
rect -1041 -114 -1025 -80
rect -991 -114 -975 -80
rect -849 -114 -833 -80
rect -799 -114 -783 -80
rect -657 -114 -641 -80
rect -607 -114 -591 -80
rect -465 -114 -449 -80
rect -415 -114 -399 -80
rect -273 -114 -257 -80
rect -223 -114 -207 -80
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect 111 -114 127 -80
rect 161 -114 177 -80
rect 303 -114 319 -80
rect 353 -114 369 -80
rect 495 -114 511 -80
rect 545 -114 561 -80
rect 687 -114 703 -80
rect 737 -114 753 -80
rect 879 -114 895 -80
rect 929 -114 945 -80
rect -1187 -182 -1153 -120
rect 1153 -182 1187 -120
rect -1187 -216 -1091 -182
rect 1091 -216 1187 -182
<< viali >>
rect -929 80 -895 114
rect -737 80 -703 114
rect -545 80 -511 114
rect -353 80 -319 114
rect -161 80 -127 114
rect 31 80 65 114
rect 223 80 257 114
rect 415 80 449 114
rect 607 80 641 114
rect 799 80 833 114
rect 991 80 1025 114
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect -1025 -114 -991 -80
rect -833 -114 -799 -80
rect -641 -114 -607 -80
rect -449 -114 -415 -80
rect -257 -114 -223 -80
rect -65 -114 -31 -80
rect 127 -114 161 -80
rect 319 -114 353 -80
rect 511 -114 545 -80
rect 703 -114 737 -80
rect 895 -114 929 -80
<< metal1 >>
rect -941 114 -883 120
rect -941 80 -929 114
rect -895 80 -883 114
rect -941 74 -883 80
rect -749 114 -691 120
rect -749 80 -737 114
rect -703 80 -691 114
rect -749 74 -691 80
rect -557 114 -499 120
rect -557 80 -545 114
rect -511 80 -499 114
rect -557 74 -499 80
rect -365 114 -307 120
rect -365 80 -353 114
rect -319 80 -307 114
rect -365 74 -307 80
rect -173 114 -115 120
rect -173 80 -161 114
rect -127 80 -115 114
rect -173 74 -115 80
rect 19 114 77 120
rect 19 80 31 114
rect 65 80 77 114
rect 19 74 77 80
rect 211 114 269 120
rect 211 80 223 114
rect 257 80 269 114
rect 211 74 269 80
rect 403 114 461 120
rect 403 80 415 114
rect 449 80 461 114
rect 403 74 461 80
rect 595 114 653 120
rect 595 80 607 114
rect 641 80 653 114
rect 595 74 653 80
rect 787 114 845 120
rect 787 80 799 114
rect 833 80 845 114
rect 787 74 845 80
rect 979 114 1037 120
rect 979 80 991 114
rect 1025 80 1037 114
rect 979 74 1037 80
rect -1079 30 -1033 42
rect -1079 -30 -1073 30
rect -1039 -30 -1033 30
rect -1079 -42 -1033 -30
rect -983 30 -937 42
rect -983 -30 -977 30
rect -943 -30 -937 30
rect -983 -42 -937 -30
rect -887 30 -841 42
rect -887 -30 -881 30
rect -847 -30 -841 30
rect -887 -42 -841 -30
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
rect 841 30 887 42
rect 841 -30 847 30
rect 881 -30 887 30
rect 841 -42 887 -30
rect 937 30 983 42
rect 937 -30 943 30
rect 977 -30 983 30
rect 937 -42 983 -30
rect 1033 30 1079 42
rect 1033 -30 1039 30
rect 1073 -30 1079 30
rect 1033 -42 1079 -30
rect -1037 -80 -979 -74
rect -1037 -114 -1025 -80
rect -991 -114 -979 -80
rect -1037 -120 -979 -114
rect -845 -80 -787 -74
rect -845 -114 -833 -80
rect -799 -114 -787 -80
rect -845 -120 -787 -114
rect -653 -80 -595 -74
rect -653 -114 -641 -80
rect -607 -114 -595 -80
rect -653 -120 -595 -114
rect -461 -80 -403 -74
rect -461 -114 -449 -80
rect -415 -114 -403 -80
rect -461 -120 -403 -114
rect -269 -80 -211 -74
rect -269 -114 -257 -80
rect -223 -114 -211 -80
rect -269 -120 -211 -114
rect -77 -80 -19 -74
rect -77 -114 -65 -80
rect -31 -114 -19 -80
rect -77 -120 -19 -114
rect 115 -80 173 -74
rect 115 -114 127 -80
rect 161 -114 173 -80
rect 115 -120 173 -114
rect 307 -80 365 -74
rect 307 -114 319 -80
rect 353 -114 365 -80
rect 307 -120 365 -114
rect 499 -80 557 -74
rect 499 -114 511 -80
rect 545 -114 557 -80
rect 499 -120 557 -114
rect 691 -80 749 -74
rect 691 -114 703 -80
rect 737 -114 749 -80
rect 691 -120 749 -114
rect 883 -80 941 -74
rect 883 -114 895 -80
rect 929 -114 941 -80
rect 883 -120 941 -114
<< properties >>
string FIXED_BBOX -1170 -199 1170 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 22 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
