magic
tech sky130A
magscale 1 2
timestamp 1695986410
<< locali >>
rect -61 170 149 1170
rect 1589 170 1765 1170
rect 46 -4 86 132
rect 1618 -4 1658 132
<< metal1 >>
rect 202 1862 254 1868
rect 202 1660 254 1666
rect 204 1170 252 1660
rect 300 1628 348 1868
rect 394 1862 446 1868
rect 394 1660 446 1666
rect 298 1622 350 1628
rect 298 1420 350 1426
rect 300 1170 348 1420
rect 396 1170 444 1660
rect 492 1628 540 1868
rect 586 1862 638 1868
rect 586 1660 638 1666
rect 490 1622 542 1628
rect 490 1420 542 1426
rect 492 1170 540 1420
rect 588 1170 636 1660
rect 684 1628 732 1868
rect 778 1862 830 1868
rect 778 1660 830 1666
rect 682 1622 734 1628
rect 682 1420 734 1426
rect 684 1170 732 1420
rect 780 1170 828 1660
rect 876 1628 924 1868
rect 970 1862 1022 1868
rect 970 1660 1022 1666
rect 874 1622 926 1628
rect 874 1420 926 1426
rect 876 1170 924 1420
rect 972 1170 1020 1660
rect 1068 1628 1116 1868
rect 1162 1862 1214 1868
rect 1162 1660 1214 1666
rect 1066 1622 1118 1628
rect 1066 1420 1118 1426
rect 1068 1170 1116 1420
rect 1164 1170 1212 1660
rect 1260 1628 1308 1868
rect 1354 1862 1406 1868
rect 1354 1660 1406 1666
rect 1258 1622 1310 1628
rect 1258 1420 1310 1426
rect 1260 1170 1308 1420
rect 1356 1170 1404 1660
rect 1452 1628 1500 1868
rect 1450 1622 1502 1628
rect 1450 1420 1502 1426
rect 1452 1170 1500 1420
rect -131 91 1835 139
<< via1 >>
rect 202 1666 254 1862
rect 394 1666 446 1862
rect 298 1426 350 1622
rect 586 1666 638 1862
rect 490 1426 542 1622
rect 778 1666 830 1862
rect 682 1426 734 1622
rect 970 1666 1022 1862
rect 874 1426 926 1622
rect 1162 1666 1214 1862
rect 1066 1426 1118 1622
rect 1354 1666 1406 1862
rect 1258 1426 1310 1622
rect 1450 1426 1502 1622
<< metal2 >>
rect 202 1862 254 1868
rect -130 1668 202 1860
rect 394 1862 446 1868
rect 254 1668 394 1860
rect 202 1660 254 1666
rect 586 1862 638 1868
rect 446 1668 586 1860
rect 394 1660 446 1666
rect 778 1862 830 1868
rect 638 1668 778 1860
rect 586 1660 638 1666
rect 970 1862 1022 1868
rect 830 1668 970 1860
rect 778 1660 830 1666
rect 1162 1862 1214 1868
rect 1022 1668 1162 1860
rect 970 1660 1022 1666
rect 1354 1862 1406 1868
rect 1214 1668 1354 1860
rect 1162 1660 1214 1666
rect 1406 1668 1842 1860
rect 1354 1660 1406 1666
rect 298 1622 350 1628
rect -130 1428 298 1620
rect 490 1622 542 1628
rect 350 1428 490 1620
rect 298 1420 350 1426
rect 682 1622 734 1628
rect 542 1428 682 1620
rect 490 1420 542 1426
rect 874 1622 926 1628
rect 734 1428 874 1620
rect 682 1420 734 1426
rect 1066 1622 1118 1628
rect 926 1428 1066 1620
rect 874 1420 926 1426
rect 1258 1622 1310 1628
rect 1118 1428 1258 1620
rect 1066 1420 1118 1426
rect 1450 1622 1502 1628
rect 1310 1428 1450 1620
rect 1258 1420 1310 1426
rect 1502 1428 1842 1620
rect 1450 1420 1502 1426
use sky130_fd_pr__nfet_01v8_YN9FL4  sky130_fd_pr__nfet_01v8_UDPJLN_0
timestamp 1695643842
transform 1 0 852 0 1 670
box -983 -710 983 710
<< labels >>
flabel locali -61 170 115 1170 0 FreeSans 240 0 0 0 vss_sw
port 0 nsew
flabel metal1 -131 91 1835 139 0 FreeSans 240 0 0 0 en_sw
port 1 nsew
<< end >>
