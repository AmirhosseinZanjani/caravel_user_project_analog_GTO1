magic
tech sky130A
magscale 1 2
timestamp 1699610342
<< pwell >>
rect 25778 29394 42564 29424
rect 25778 28864 42566 29394
rect 39838 24242 41330 28864
<< locali >>
rect 6414 291908 8494 291994
rect 6414 291560 6492 291908
rect 8288 291560 8494 291908
rect 6414 20004 8494 291560
rect 49366 58822 67588 58862
rect 24812 58556 91822 58822
rect 24812 57078 50752 58556
rect 61688 57078 91822 58556
rect 24812 56840 91822 57078
rect 24816 49868 30784 56840
rect 24816 33856 30792 49868
rect 57284 44892 59236 56840
rect 57308 44476 57818 44892
rect 89738 44358 91690 56840
rect 30458 33848 30792 33856
rect 24812 31140 30754 31160
rect 24796 31044 30754 31140
rect 24796 29424 30748 31044
rect 24796 29394 42564 29424
rect 24796 29360 42566 29394
rect 24796 28906 24854 29360
rect 25320 28906 42566 29360
rect 24796 28864 42566 28906
rect 24796 28856 30748 28864
rect 39838 24242 41330 28864
rect 6414 19998 20564 20004
rect 6414 19996 33806 19998
rect 6414 19872 36062 19996
rect 6414 19412 34304 19872
rect 35416 19412 36062 19872
rect 6414 19352 36062 19412
rect 6414 19350 20564 19352
rect 32376 19350 36062 19352
<< viali >>
rect 6492 291560 8288 291908
rect 50752 57078 61688 58556
rect 24854 28906 25320 29360
rect 34304 19412 35416 19872
<< metal1 >>
rect 38932 696022 40588 696178
rect 38932 692550 38950 696022
rect 40550 692550 40588 696022
rect 12450 685220 14128 685300
rect 12440 680274 12450 685220
rect 14082 683684 14128 685220
rect 14082 680274 14138 683684
rect 12450 556104 14138 680274
rect 38932 680262 40588 692550
rect 12450 549442 14122 556104
rect 6390 291210 6400 291992
rect 8504 291210 8514 291992
rect 12450 32152 14138 549442
rect 38932 32168 40620 680262
rect 72242 378424 75630 378428
rect 72234 377956 72244 378424
rect 75638 377956 75648 378424
rect 50042 56728 50052 59732
rect 62538 56728 62548 59732
rect 72242 47074 75630 377956
rect 72222 44890 72232 46422
rect 75674 44890 75684 46422
rect 22164 32152 26952 32154
rect 12450 31982 26952 32152
rect 28620 31982 40620 32168
rect 20262 31976 26952 31982
rect 22164 31974 26952 31976
rect 28628 31980 33416 31982
rect 26806 31738 26944 31974
rect 28628 31744 28766 31980
rect 38932 31970 40620 31982
rect 27312 30452 27480 31262
rect 27312 30368 27482 30452
rect 22860 29454 25714 29870
rect 22814 29440 25756 29454
rect 22814 28906 22882 29440
rect 23962 29360 25756 29440
rect 23962 28906 24854 29360
rect 25320 28906 25756 29360
rect 27314 29032 27482 30368
rect 28084 29032 28250 31256
rect 27314 28940 28252 29032
rect 22814 28860 25756 28906
rect 22860 27798 25714 28860
rect 27318 28802 28252 28940
rect 27312 7324 28254 28802
rect 73720 22378 73730 23234
rect 75120 22378 75130 23234
rect 36002 19986 36820 20016
rect 34268 19872 36820 19986
rect 34268 19412 34304 19872
rect 35416 19412 36820 19872
rect 34268 19360 36820 19412
rect 44164 19360 94568 19986
rect 36002 16300 36820 19360
rect 73734 16300 75152 19360
rect 36002 15348 75152 16300
rect 36002 15314 36820 15348
rect 73734 15316 75152 15348
rect 578740 7324 578750 7342
rect 27312 3046 578750 7324
rect 579820 3046 579830 7342
<< via1 >>
rect 38950 692550 40550 696022
rect 12450 680274 14082 685220
rect 6400 291908 8504 291992
rect 6400 291560 6492 291908
rect 6492 291560 8288 291908
rect 8288 291560 8504 291908
rect 6400 291210 8504 291560
rect 72244 377956 75638 378424
rect 50052 58556 62538 59732
rect 50052 57078 50752 58556
rect 50752 57078 61688 58556
rect 61688 57078 62538 58556
rect 50052 56728 62538 57078
rect 72232 44890 75674 46422
rect 22882 28906 23962 29440
rect 73730 22378 75120 23234
rect 578750 3046 579820 7342
<< metal2 >>
rect 38940 696022 40550 696032
rect 38940 692540 40550 692550
rect 12450 685220 14082 685230
rect 12450 680264 14082 680274
rect 67540 580218 73832 580228
rect 67540 574370 73832 574380
rect 67666 490684 73818 574370
rect 120256 502524 125154 502534
rect 103538 500856 120256 501886
rect 103510 498372 120256 500856
rect 67666 463324 73816 490684
rect 44418 461296 73816 463324
rect 44422 335208 45414 461296
rect 67666 460568 73816 461296
rect 72244 378424 75638 378434
rect 72244 377946 75638 377956
rect 72760 335214 75250 335224
rect 44420 335096 45414 335208
rect 72758 335096 72760 335208
rect 6400 291992 8504 292002
rect 6400 291200 8504 291210
rect 3674 248982 5612 248992
rect 3672 248656 3674 248970
rect 3672 7050 5612 248656
rect 21552 29768 24406 29870
rect 21552 28854 21622 29768
rect 23968 28854 24406 29768
rect 21552 27914 21648 28854
rect 23956 27914 24406 28854
rect 26214 28624 26352 31048
rect 21552 27798 24406 27914
rect 26210 28278 26352 28624
rect 44422 28310 45414 335096
rect 75250 335024 75252 335212
rect 72760 335014 75252 335024
rect 72768 334352 75252 335014
rect 50052 59732 62538 59742
rect 50052 56718 62538 56728
rect 72768 46432 75262 334352
rect 72232 46422 75674 46432
rect 72232 44880 75674 44890
rect 51678 28310 58914 28314
rect 26210 23898 26350 28278
rect 44422 28072 58914 28310
rect 103510 28248 104514 498372
rect 120256 498148 125154 498158
rect 85432 28094 104514 28248
rect 103510 28076 104514 28094
rect 44422 28066 52902 28072
rect 26210 23666 26352 23898
rect 26214 8746 26352 23666
rect 73730 23236 75120 23244
rect 73716 23234 75348 23236
rect 73716 22378 73730 23234
rect 75120 22378 75348 23234
rect 73716 16548 75348 22378
rect 73716 13484 75394 16548
rect 26214 8626 26352 8636
rect 73762 7100 75394 13484
rect 23222 7052 75394 7100
rect 9760 7050 75394 7052
rect 3672 6796 75394 7050
rect 578750 7342 579820 7352
rect 3672 4664 75362 6796
rect 3672 4568 24768 4664
rect 3672 4566 19600 4568
rect 3672 4562 5612 4566
rect 578750 3036 579820 3046
rect 579704 -800 579820 3036
<< via2 >>
rect 38940 692550 38950 696022
rect 38950 692550 40550 696022
rect 12450 680274 14082 685220
rect 67540 574380 73832 580218
rect 72244 377956 75638 378424
rect 6400 291210 8504 291992
rect 3674 248656 5612 248982
rect 21622 29440 23968 29768
rect 21622 28906 22882 29440
rect 22882 28906 23962 29440
rect 23962 28906 23968 29440
rect 21622 28854 23968 28906
rect 21648 27914 23956 28854
rect 72760 335024 75250 335214
rect 50052 56728 62538 59732
rect 120256 498158 125154 502524
rect 26214 8636 26352 8746
<< metal3 >>
rect 16168 696218 21162 704916
rect 16168 696140 40628 696218
rect 16208 696022 40628 696140
rect 16208 692550 38940 696022
rect 40550 692550 40628 696022
rect 38930 692545 40560 692550
rect -800 685220 14136 685278
rect -800 680274 12450 685220
rect 14082 680274 14136 685220
rect -800 680242 14136 680274
rect 68190 580223 73194 702712
rect 120202 695584 125188 703972
rect 67530 580218 73842 580223
rect 67530 574380 67540 580218
rect 73832 574380 73842 580218
rect 67530 574375 73842 574380
rect -1600 562412 23964 564306
rect -1600 560772 15446 562412
rect 20410 560772 23964 562412
rect -1600 559442 23964 560772
rect -800 549442 866 554278
rect 120202 502524 125190 695584
rect 120202 500158 120256 502524
rect 120246 498158 120256 500158
rect 125154 500158 125190 502524
rect 125154 498158 125164 500158
rect 120246 498153 125164 498158
rect -800 378428 71758 378432
rect 72234 378428 75648 378429
rect -800 378424 75648 378428
rect -800 378318 72244 378424
rect 72234 377956 72244 378318
rect 75638 377956 75648 378424
rect 72234 377951 75648 377956
rect 72750 335214 75260 335219
rect 72750 335208 72760 335214
rect -800 335096 72760 335208
rect 72750 335024 72760 335096
rect 75250 335024 75260 335214
rect 72750 335019 75260 335024
rect 6390 291992 8514 291997
rect -800 291874 6400 291992
rect 6390 291210 6400 291874
rect 8504 291210 8514 291992
rect 6390 291205 8514 291210
rect 3664 248982 5622 248987
rect -800 248964 2748 248966
rect 3664 248964 3674 248982
rect -800 248852 3674 248964
rect 3664 248656 3674 248852
rect 5612 248656 5622 248982
rect 3664 248651 5622 248656
rect -800 209622 11482 209690
rect -800 209462 44374 209622
rect -800 204888 62556 209462
rect 11542 64458 23914 65596
rect 11542 55812 12568 64458
rect 23264 55812 23914 64458
rect 50184 59737 62556 204888
rect 50042 59732 62556 59737
rect 50042 56728 50052 59732
rect 62538 56728 62556 59732
rect 50042 56723 62548 56728
rect 11542 30152 23914 55812
rect 107686 35204 108194 35254
rect 38330 34876 55606 35168
rect 11542 29768 23986 30152
rect 11542 28854 21622 29768
rect 23968 28854 23986 29768
rect 11542 27914 21648 28854
rect 23956 28176 23986 28854
rect 23956 27914 23966 28176
rect 11542 27909 23966 27914
rect 11542 27802 23914 27909
rect 29256 27370 29390 31048
rect 29256 26752 29392 27370
rect 29256 26748 29394 26752
rect 29256 26066 29396 26748
rect 38330 26066 39256 34876
rect 91070 34792 108194 35204
rect 29176 24796 39282 26066
rect 29256 21066 29394 24796
rect 29254 20432 29394 21066
rect 29254 17090 29392 20432
rect 29254 17086 29394 17090
rect 29256 16162 29394 17086
rect 29252 13110 29394 16162
rect -800 12294 27254 12296
rect -800 12288 27914 12294
rect 29252 12288 29390 13110
rect -800 12182 29400 12288
rect 107686 11800 108194 34792
rect -800 8746 12044 8748
rect 26204 8746 26362 8751
rect -800 8636 26214 8746
rect 26352 8730 26362 8746
rect 107686 8730 108162 11800
rect 26352 8636 108162 8730
rect 26204 8631 26362 8636
rect 107686 8596 108162 8636
<< via3 >>
rect 15446 560772 20410 562412
rect 12568 55812 23264 64458
<< metal4 >>
rect 11658 562412 23922 564264
rect 11658 560772 15446 562412
rect 20410 560772 23922 562412
rect 11658 383278 23922 560772
rect 11658 64458 24170 383278
rect 11658 56038 12568 64458
rect 12567 55812 12568 56038
rect 23264 56038 24170 64458
rect 23264 55812 23265 56038
rect 12567 55811 23265 55812
use integrator  integrator_0
timestamp 1699562254
transform 1 0 41328 0 1 24550
box -66 -5190 66178 23186
use Quantizer  Quantizer_0
timestamp 1699568647
transform 1 0 24915 0 1 31120
box -137 -142 5874 3158
<< end >>
