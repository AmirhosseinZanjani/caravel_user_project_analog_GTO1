magic
tech sky130A
magscale 1 2
timestamp 1696338270
use capbank  capbank_0
timestamp 1696325208
transform 1 0 8083 0 1 -10120
box -4432 -9317 8974 20462
use osc_total  osc_total_0
timestamp 1696337502
transform 1 0 0 0 1 0
box -3210 -7260 23916 29082
use uwb_inductor  uwb_inductor_0
timestamp 1695396033
transform 1 0 10352 0 1 12240
box -9750 -1500 9750 18750
<< end >>
