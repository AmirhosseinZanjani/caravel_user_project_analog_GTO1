magic
tech sky130A
magscale 1 2
timestamp 1695991705
<< via2 >>
rect 1836 17956 2146 18148
rect 2396 17716 2706 17908
rect 1836 11638 2146 11830
rect 2396 11398 2706 11590
<< metal3 >>
rect 1806 18166 2176 18196
rect 1806 17640 1836 18166
rect 2146 17640 2176 18166
rect 1806 17610 2176 17640
rect 2366 18166 2736 18196
rect 2366 17640 2396 18166
rect 2706 17640 2736 18166
rect 2366 17610 2736 17640
rect 1806 11848 2176 11878
rect 1806 11322 1836 11848
rect 2146 11322 2176 11848
rect 1806 11292 2176 11322
rect 2366 11848 2736 11878
rect 2366 11322 2396 11848
rect 2706 11322 2736 11848
rect 2366 11292 2736 11322
<< via3 >>
rect 1836 18148 2146 18166
rect 1836 17956 2146 18148
rect 1836 17640 2146 17956
rect 2396 17908 2706 18166
rect 2396 17716 2706 17908
rect 2396 17640 2706 17716
rect 1836 11830 2146 11848
rect 1836 11638 2146 11830
rect 1836 11322 2146 11638
rect 2396 11590 2706 11848
rect 2396 11398 2706 11590
rect 2396 11322 2706 11398
<< metal4 >>
rect 2366 19706 2736 19710
rect -3844 19680 2176 19706
rect -3844 19370 -3430 19680
rect -2490 19370 2176 19680
rect -3844 19336 2176 19370
rect -3844 18490 1176 18524
rect -3844 17900 -1948 18490
rect -1208 17900 1176 18490
rect -3844 17874 1176 17900
rect 1806 18166 2176 19336
rect 1806 17640 1836 18166
rect 2146 17640 2176 18166
rect 1806 17610 2176 17640
rect 2366 19680 8386 19706
rect 2366 19370 7030 19680
rect 7970 19370 8386 19680
rect 2366 19336 8386 19370
rect 2366 18166 2736 19336
rect 2366 17640 2396 18166
rect 2706 17640 2736 18166
rect 3366 18490 8386 18524
rect 3366 17900 5750 18490
rect 6490 17900 8386 18490
rect 3366 17874 8386 17900
rect 2366 17610 2736 17640
rect -3844 17030 1176 17062
rect -3844 16440 -3430 17030
rect -2490 16440 1176 17030
rect -3844 16412 1176 16440
rect 3366 17030 8386 17062
rect 3366 16440 7030 17030
rect 7970 16440 8386 17030
rect 3366 16412 8386 16440
rect -3844 15570 1176 15600
rect -3844 14980 -1948 15570
rect -1208 14980 1176 15570
rect -3844 14950 1176 14980
rect 3366 15570 8386 15600
rect 3366 14980 5750 15570
rect 6490 14980 8386 15570
rect 3366 14950 8386 14980
rect -3844 14110 1176 14138
rect -3844 13800 -3430 14110
rect -2490 13800 1176 14110
rect -3844 13768 1176 13800
rect 3366 14110 8386 14138
rect 3366 13800 7030 14110
rect 7970 13800 8386 14110
rect 3366 13768 8386 13800
rect -3844 13360 2176 13388
rect -3844 13050 -3428 13360
rect -2488 13050 2176 13360
rect -3844 13018 2176 13050
rect -3844 12176 1176 12206
rect -3844 11586 -1948 12176
rect -1208 11586 1176 12176
rect -3844 11556 1176 11586
rect 1806 11848 2176 13018
rect 1806 11322 1836 11848
rect 2146 11322 2176 11848
rect 1806 11292 2176 11322
rect 2366 13360 8386 13388
rect 2366 13050 7030 13360
rect 7970 13050 8386 13360
rect 2366 13018 8386 13050
rect 2366 11848 2736 13018
rect 2366 11322 2396 11848
rect 2706 11322 2736 11848
rect 3366 12176 8386 12206
rect 3366 11586 5750 12176
rect 6490 11586 8386 12176
rect 3366 11556 8386 11586
rect 2366 11292 2736 11322
rect -3844 10716 1176 10746
rect -3844 10126 -3428 10716
rect -2488 10126 1176 10716
rect -3844 10096 1176 10126
rect 3366 10716 8386 10746
rect 3366 10126 7030 10716
rect 7970 10126 8386 10716
rect 3366 10096 8386 10126
rect -3844 9256 1176 9286
rect -3844 8666 -1948 9256
rect -1208 8666 1176 9256
rect -3844 8636 1176 8666
rect 3366 9256 8386 9286
rect 3366 8666 5750 9256
rect 6490 8666 8386 9256
rect 3366 8636 8386 8666
rect -3844 7788 1176 7820
rect -3844 7478 -3428 7788
rect -2488 7478 1176 7788
rect -3844 7450 1176 7478
rect 3366 7790 8386 7820
rect 3366 7480 7030 7790
rect 7970 7480 8386 7790
rect 3366 7450 8386 7480
<< via4 >>
rect -3430 19370 -2490 19680
rect -1948 17900 -1208 18490
rect 7030 19370 7970 19680
rect 5750 17900 6490 18490
rect -3430 16440 -2490 17030
rect 7030 16440 7970 17030
rect -1948 14980 -1208 15570
rect 5750 14980 6490 15570
rect -3430 13800 -2490 14110
rect 7030 13800 7970 14110
rect -3428 13050 -2488 13360
rect -1948 11586 -1208 12176
rect 7030 13050 7970 13360
rect 5750 11586 6490 12176
rect -3428 10126 -2488 10716
rect 7030 10126 7970 10716
rect -1948 8666 -1208 9256
rect 5750 8666 6490 9256
rect -3428 7478 -2488 7788
rect 7030 7480 7970 7790
<< metal5 >>
rect -3457 19680 -2457 19706
rect -3457 19370 -3430 19680
rect -2490 19370 -2457 19680
rect -3457 17030 -2457 19370
rect -1457 18530 -457 20462
rect -1980 18490 -457 18530
rect -1980 17900 -1948 18490
rect -1208 17900 -457 18490
rect -1980 17870 -457 17900
rect -3457 16440 -3430 17030
rect -2490 16440 -2457 17030
rect -3457 14110 -2457 16440
rect -1457 15600 -457 17870
rect -1980 15570 -457 15600
rect -1980 14980 -1948 15570
rect -1208 14980 -457 15570
rect -1980 14950 -457 14980
rect -3457 13800 -3430 14110
rect -2490 13800 -2457 14110
rect -3457 13768 -2457 13800
rect -3457 13360 -2457 13388
rect -3457 13050 -3428 13360
rect -2488 13050 -2457 13360
rect -3457 10716 -2457 13050
rect -1457 12206 -457 14950
rect -1978 12176 -457 12206
rect -1978 11586 -1948 12176
rect -1208 11586 -457 12176
rect -1978 11556 -457 11586
rect -3457 10126 -3428 10716
rect -2488 10126 -2457 10716
rect -3457 7788 -2457 10126
rect -1457 9286 -457 11556
rect -1978 9256 -457 9286
rect -1978 8666 -1948 9256
rect -1208 8666 -457 9256
rect -1978 8636 -457 8666
rect -3457 7478 -3428 7788
rect -2488 7478 -2457 7788
rect -3457 7450 -2457 7478
rect -1457 -2738 -457 8636
rect 4999 18530 6000 20462
rect 6999 19680 8000 19706
rect 6999 19370 7030 19680
rect 7970 19370 8000 19680
rect 4999 18490 6520 18530
rect 4999 17900 5750 18490
rect 6490 17900 6520 18490
rect 4999 17870 6520 17900
rect 4999 15600 6000 17870
rect 6999 17030 8000 19370
rect 6999 16440 7030 17030
rect 7970 16440 8000 17030
rect 4999 15570 6520 15600
rect 4999 14980 5750 15570
rect 6490 14980 6520 15570
rect 4999 14950 6520 14980
rect 4999 12206 6000 14950
rect 6999 14110 8000 16440
rect 6999 13800 7030 14110
rect 7970 13800 8000 14110
rect 6999 13768 8000 13800
rect 6999 13360 8000 13388
rect 6999 13050 7030 13360
rect 7970 13050 8000 13360
rect 4999 12176 6520 12206
rect 4999 11586 5750 12176
rect 6490 11586 6520 12176
rect 4999 11556 6520 11586
rect 4999 9286 6000 11556
rect 6999 10716 8000 13050
rect 6999 10126 7030 10716
rect 7970 10126 8000 10716
rect 4999 9256 6520 9286
rect 4999 8666 5750 9256
rect 6490 8666 6520 9256
rect 4999 8636 6520 8666
rect 4999 -2738 6000 8636
rect 6999 7790 8000 10126
rect 6999 7480 7030 7790
rect 7970 7480 8000 7790
rect 6999 7450 8000 7480
use capbank_1  capbank_1_0
timestamp 1695986410
transform 1 0 1288 0 -1 -816
box -1292 0 3258 1908
use capbank_2  capbank_2_0
timestamp 1695986410
transform 1 0 1288 0 -1 1092
box -2572 0 4538 1908
use capbank_4  capbank_4_0
timestamp 1695986410
transform 1 0 1288 0 -1 4216
box -2572 0 4538 2834
use capbank_8  capbank_8_1
timestamp 1695986410
transform 1 0 1288 0 -1 7340
box -5132 0 7098 2834
use capbank_16  capbank_16_0
timestamp 1695986410
transform 1 0 1288 0 -1 19616
box -5132 0 7098 5758
use capbank_16  capbank_16_1
timestamp 1695986410
transform 1 0 1288 0 -1 13298
box -5132 0 7098 5758
use uwb_inductor  uwb_inductor_0
timestamp 1695396033
transform 1 0 2271 0 1 22362
box -9750 -1500 9750 18750
<< end >>
