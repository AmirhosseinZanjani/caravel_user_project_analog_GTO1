magic
tech sky130A
magscale 1 2
timestamp 1697034114
<< nwell >>
rect -11321 -319 11321 319
<< pmos >>
rect -11125 -100 -10325 100
rect -10267 -100 -9467 100
rect -9409 -100 -8609 100
rect -8551 -100 -7751 100
rect -7693 -100 -6893 100
rect -6835 -100 -6035 100
rect -5977 -100 -5177 100
rect -5119 -100 -4319 100
rect -4261 -100 -3461 100
rect -3403 -100 -2603 100
rect -2545 -100 -1745 100
rect -1687 -100 -887 100
rect -829 -100 -29 100
rect 29 -100 829 100
rect 887 -100 1687 100
rect 1745 -100 2545 100
rect 2603 -100 3403 100
rect 3461 -100 4261 100
rect 4319 -100 5119 100
rect 5177 -100 5977 100
rect 6035 -100 6835 100
rect 6893 -100 7693 100
rect 7751 -100 8551 100
rect 8609 -100 9409 100
rect 9467 -100 10267 100
rect 10325 -100 11125 100
<< pdiff >>
rect -11183 88 -11125 100
rect -11183 -88 -11171 88
rect -11137 -88 -11125 88
rect -11183 -100 -11125 -88
rect -10325 88 -10267 100
rect -10325 -88 -10313 88
rect -10279 -88 -10267 88
rect -10325 -100 -10267 -88
rect -9467 88 -9409 100
rect -9467 -88 -9455 88
rect -9421 -88 -9409 88
rect -9467 -100 -9409 -88
rect -8609 88 -8551 100
rect -8609 -88 -8597 88
rect -8563 -88 -8551 88
rect -8609 -100 -8551 -88
rect -7751 88 -7693 100
rect -7751 -88 -7739 88
rect -7705 -88 -7693 88
rect -7751 -100 -7693 -88
rect -6893 88 -6835 100
rect -6893 -88 -6881 88
rect -6847 -88 -6835 88
rect -6893 -100 -6835 -88
rect -6035 88 -5977 100
rect -6035 -88 -6023 88
rect -5989 -88 -5977 88
rect -6035 -100 -5977 -88
rect -5177 88 -5119 100
rect -5177 -88 -5165 88
rect -5131 -88 -5119 88
rect -5177 -100 -5119 -88
rect -4319 88 -4261 100
rect -4319 -88 -4307 88
rect -4273 -88 -4261 88
rect -4319 -100 -4261 -88
rect -3461 88 -3403 100
rect -3461 -88 -3449 88
rect -3415 -88 -3403 88
rect -3461 -100 -3403 -88
rect -2603 88 -2545 100
rect -2603 -88 -2591 88
rect -2557 -88 -2545 88
rect -2603 -100 -2545 -88
rect -1745 88 -1687 100
rect -1745 -88 -1733 88
rect -1699 -88 -1687 88
rect -1745 -100 -1687 -88
rect -887 88 -829 100
rect -887 -88 -875 88
rect -841 -88 -829 88
rect -887 -100 -829 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 829 88 887 100
rect 829 -88 841 88
rect 875 -88 887 88
rect 829 -100 887 -88
rect 1687 88 1745 100
rect 1687 -88 1699 88
rect 1733 -88 1745 88
rect 1687 -100 1745 -88
rect 2545 88 2603 100
rect 2545 -88 2557 88
rect 2591 -88 2603 88
rect 2545 -100 2603 -88
rect 3403 88 3461 100
rect 3403 -88 3415 88
rect 3449 -88 3461 88
rect 3403 -100 3461 -88
rect 4261 88 4319 100
rect 4261 -88 4273 88
rect 4307 -88 4319 88
rect 4261 -100 4319 -88
rect 5119 88 5177 100
rect 5119 -88 5131 88
rect 5165 -88 5177 88
rect 5119 -100 5177 -88
rect 5977 88 6035 100
rect 5977 -88 5989 88
rect 6023 -88 6035 88
rect 5977 -100 6035 -88
rect 6835 88 6893 100
rect 6835 -88 6847 88
rect 6881 -88 6893 88
rect 6835 -100 6893 -88
rect 7693 88 7751 100
rect 7693 -88 7705 88
rect 7739 -88 7751 88
rect 7693 -100 7751 -88
rect 8551 88 8609 100
rect 8551 -88 8563 88
rect 8597 -88 8609 88
rect 8551 -100 8609 -88
rect 9409 88 9467 100
rect 9409 -88 9421 88
rect 9455 -88 9467 88
rect 9409 -100 9467 -88
rect 10267 88 10325 100
rect 10267 -88 10279 88
rect 10313 -88 10325 88
rect 10267 -100 10325 -88
rect 11125 88 11183 100
rect 11125 -88 11137 88
rect 11171 -88 11183 88
rect 11125 -100 11183 -88
<< pdiffc >>
rect -11171 -88 -11137 88
rect -10313 -88 -10279 88
rect -9455 -88 -9421 88
rect -8597 -88 -8563 88
rect -7739 -88 -7705 88
rect -6881 -88 -6847 88
rect -6023 -88 -5989 88
rect -5165 -88 -5131 88
rect -4307 -88 -4273 88
rect -3449 -88 -3415 88
rect -2591 -88 -2557 88
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect 2557 -88 2591 88
rect 3415 -88 3449 88
rect 4273 -88 4307 88
rect 5131 -88 5165 88
rect 5989 -88 6023 88
rect 6847 -88 6881 88
rect 7705 -88 7739 88
rect 8563 -88 8597 88
rect 9421 -88 9455 88
rect 10279 -88 10313 88
rect 11137 -88 11171 88
<< nsubdiff >>
rect -11285 249 -11189 283
rect 11189 249 11285 283
rect -11285 187 -11251 249
rect 11251 187 11285 249
rect -11285 -249 -11251 -187
rect 11251 -249 11285 -187
rect -11285 -283 -11189 -249
rect 11189 -283 11285 -249
<< nsubdiffcont >>
rect -11189 249 11189 283
rect -11285 -187 -11251 187
rect 11251 -187 11285 187
rect -11189 -283 11189 -249
<< poly >>
rect -11125 181 -10325 197
rect -11125 147 -11109 181
rect -10341 147 -10325 181
rect -11125 100 -10325 147
rect -10267 181 -9467 197
rect -10267 147 -10251 181
rect -9483 147 -9467 181
rect -10267 100 -9467 147
rect -9409 181 -8609 197
rect -9409 147 -9393 181
rect -8625 147 -8609 181
rect -9409 100 -8609 147
rect -8551 181 -7751 197
rect -8551 147 -8535 181
rect -7767 147 -7751 181
rect -8551 100 -7751 147
rect -7693 181 -6893 197
rect -7693 147 -7677 181
rect -6909 147 -6893 181
rect -7693 100 -6893 147
rect -6835 181 -6035 197
rect -6835 147 -6819 181
rect -6051 147 -6035 181
rect -6835 100 -6035 147
rect -5977 181 -5177 197
rect -5977 147 -5961 181
rect -5193 147 -5177 181
rect -5977 100 -5177 147
rect -5119 181 -4319 197
rect -5119 147 -5103 181
rect -4335 147 -4319 181
rect -5119 100 -4319 147
rect -4261 181 -3461 197
rect -4261 147 -4245 181
rect -3477 147 -3461 181
rect -4261 100 -3461 147
rect -3403 181 -2603 197
rect -3403 147 -3387 181
rect -2619 147 -2603 181
rect -3403 100 -2603 147
rect -2545 181 -1745 197
rect -2545 147 -2529 181
rect -1761 147 -1745 181
rect -2545 100 -1745 147
rect -1687 181 -887 197
rect -1687 147 -1671 181
rect -903 147 -887 181
rect -1687 100 -887 147
rect -829 181 -29 197
rect -829 147 -813 181
rect -45 147 -29 181
rect -829 100 -29 147
rect 29 181 829 197
rect 29 147 45 181
rect 813 147 829 181
rect 29 100 829 147
rect 887 181 1687 197
rect 887 147 903 181
rect 1671 147 1687 181
rect 887 100 1687 147
rect 1745 181 2545 197
rect 1745 147 1761 181
rect 2529 147 2545 181
rect 1745 100 2545 147
rect 2603 181 3403 197
rect 2603 147 2619 181
rect 3387 147 3403 181
rect 2603 100 3403 147
rect 3461 181 4261 197
rect 3461 147 3477 181
rect 4245 147 4261 181
rect 3461 100 4261 147
rect 4319 181 5119 197
rect 4319 147 4335 181
rect 5103 147 5119 181
rect 4319 100 5119 147
rect 5177 181 5977 197
rect 5177 147 5193 181
rect 5961 147 5977 181
rect 5177 100 5977 147
rect 6035 181 6835 197
rect 6035 147 6051 181
rect 6819 147 6835 181
rect 6035 100 6835 147
rect 6893 181 7693 197
rect 6893 147 6909 181
rect 7677 147 7693 181
rect 6893 100 7693 147
rect 7751 181 8551 197
rect 7751 147 7767 181
rect 8535 147 8551 181
rect 7751 100 8551 147
rect 8609 181 9409 197
rect 8609 147 8625 181
rect 9393 147 9409 181
rect 8609 100 9409 147
rect 9467 181 10267 197
rect 9467 147 9483 181
rect 10251 147 10267 181
rect 9467 100 10267 147
rect 10325 181 11125 197
rect 10325 147 10341 181
rect 11109 147 11125 181
rect 10325 100 11125 147
rect -11125 -147 -10325 -100
rect -11125 -181 -11109 -147
rect -10341 -181 -10325 -147
rect -11125 -197 -10325 -181
rect -10267 -147 -9467 -100
rect -10267 -181 -10251 -147
rect -9483 -181 -9467 -147
rect -10267 -197 -9467 -181
rect -9409 -147 -8609 -100
rect -9409 -181 -9393 -147
rect -8625 -181 -8609 -147
rect -9409 -197 -8609 -181
rect -8551 -147 -7751 -100
rect -8551 -181 -8535 -147
rect -7767 -181 -7751 -147
rect -8551 -197 -7751 -181
rect -7693 -147 -6893 -100
rect -7693 -181 -7677 -147
rect -6909 -181 -6893 -147
rect -7693 -197 -6893 -181
rect -6835 -147 -6035 -100
rect -6835 -181 -6819 -147
rect -6051 -181 -6035 -147
rect -6835 -197 -6035 -181
rect -5977 -147 -5177 -100
rect -5977 -181 -5961 -147
rect -5193 -181 -5177 -147
rect -5977 -197 -5177 -181
rect -5119 -147 -4319 -100
rect -5119 -181 -5103 -147
rect -4335 -181 -4319 -147
rect -5119 -197 -4319 -181
rect -4261 -147 -3461 -100
rect -4261 -181 -4245 -147
rect -3477 -181 -3461 -147
rect -4261 -197 -3461 -181
rect -3403 -147 -2603 -100
rect -3403 -181 -3387 -147
rect -2619 -181 -2603 -147
rect -3403 -197 -2603 -181
rect -2545 -147 -1745 -100
rect -2545 -181 -2529 -147
rect -1761 -181 -1745 -147
rect -2545 -197 -1745 -181
rect -1687 -147 -887 -100
rect -1687 -181 -1671 -147
rect -903 -181 -887 -147
rect -1687 -197 -887 -181
rect -829 -147 -29 -100
rect -829 -181 -813 -147
rect -45 -181 -29 -147
rect -829 -197 -29 -181
rect 29 -147 829 -100
rect 29 -181 45 -147
rect 813 -181 829 -147
rect 29 -197 829 -181
rect 887 -147 1687 -100
rect 887 -181 903 -147
rect 1671 -181 1687 -147
rect 887 -197 1687 -181
rect 1745 -147 2545 -100
rect 1745 -181 1761 -147
rect 2529 -181 2545 -147
rect 1745 -197 2545 -181
rect 2603 -147 3403 -100
rect 2603 -181 2619 -147
rect 3387 -181 3403 -147
rect 2603 -197 3403 -181
rect 3461 -147 4261 -100
rect 3461 -181 3477 -147
rect 4245 -181 4261 -147
rect 3461 -197 4261 -181
rect 4319 -147 5119 -100
rect 4319 -181 4335 -147
rect 5103 -181 5119 -147
rect 4319 -197 5119 -181
rect 5177 -147 5977 -100
rect 5177 -181 5193 -147
rect 5961 -181 5977 -147
rect 5177 -197 5977 -181
rect 6035 -147 6835 -100
rect 6035 -181 6051 -147
rect 6819 -181 6835 -147
rect 6035 -197 6835 -181
rect 6893 -147 7693 -100
rect 6893 -181 6909 -147
rect 7677 -181 7693 -147
rect 6893 -197 7693 -181
rect 7751 -147 8551 -100
rect 7751 -181 7767 -147
rect 8535 -181 8551 -147
rect 7751 -197 8551 -181
rect 8609 -147 9409 -100
rect 8609 -181 8625 -147
rect 9393 -181 9409 -147
rect 8609 -197 9409 -181
rect 9467 -147 10267 -100
rect 9467 -181 9483 -147
rect 10251 -181 10267 -147
rect 9467 -197 10267 -181
rect 10325 -147 11125 -100
rect 10325 -181 10341 -147
rect 11109 -181 11125 -147
rect 10325 -197 11125 -181
<< polycont >>
rect -11109 147 -10341 181
rect -10251 147 -9483 181
rect -9393 147 -8625 181
rect -8535 147 -7767 181
rect -7677 147 -6909 181
rect -6819 147 -6051 181
rect -5961 147 -5193 181
rect -5103 147 -4335 181
rect -4245 147 -3477 181
rect -3387 147 -2619 181
rect -2529 147 -1761 181
rect -1671 147 -903 181
rect -813 147 -45 181
rect 45 147 813 181
rect 903 147 1671 181
rect 1761 147 2529 181
rect 2619 147 3387 181
rect 3477 147 4245 181
rect 4335 147 5103 181
rect 5193 147 5961 181
rect 6051 147 6819 181
rect 6909 147 7677 181
rect 7767 147 8535 181
rect 8625 147 9393 181
rect 9483 147 10251 181
rect 10341 147 11109 181
rect -11109 -181 -10341 -147
rect -10251 -181 -9483 -147
rect -9393 -181 -8625 -147
rect -8535 -181 -7767 -147
rect -7677 -181 -6909 -147
rect -6819 -181 -6051 -147
rect -5961 -181 -5193 -147
rect -5103 -181 -4335 -147
rect -4245 -181 -3477 -147
rect -3387 -181 -2619 -147
rect -2529 -181 -1761 -147
rect -1671 -181 -903 -147
rect -813 -181 -45 -147
rect 45 -181 813 -147
rect 903 -181 1671 -147
rect 1761 -181 2529 -147
rect 2619 -181 3387 -147
rect 3477 -181 4245 -147
rect 4335 -181 5103 -147
rect 5193 -181 5961 -147
rect 6051 -181 6819 -147
rect 6909 -181 7677 -147
rect 7767 -181 8535 -147
rect 8625 -181 9393 -147
rect 9483 -181 10251 -147
rect 10341 -181 11109 -147
<< locali >>
rect -11285 249 -11189 283
rect 11189 249 11285 283
rect -11285 187 -11251 249
rect 11251 187 11285 249
rect -11125 147 -11109 181
rect -10341 147 -10325 181
rect -10267 147 -10251 181
rect -9483 147 -9467 181
rect -9409 147 -9393 181
rect -8625 147 -8609 181
rect -8551 147 -8535 181
rect -7767 147 -7751 181
rect -7693 147 -7677 181
rect -6909 147 -6893 181
rect -6835 147 -6819 181
rect -6051 147 -6035 181
rect -5977 147 -5961 181
rect -5193 147 -5177 181
rect -5119 147 -5103 181
rect -4335 147 -4319 181
rect -4261 147 -4245 181
rect -3477 147 -3461 181
rect -3403 147 -3387 181
rect -2619 147 -2603 181
rect -2545 147 -2529 181
rect -1761 147 -1745 181
rect -1687 147 -1671 181
rect -903 147 -887 181
rect -829 147 -813 181
rect -45 147 -29 181
rect 29 147 45 181
rect 813 147 829 181
rect 887 147 903 181
rect 1671 147 1687 181
rect 1745 147 1761 181
rect 2529 147 2545 181
rect 2603 147 2619 181
rect 3387 147 3403 181
rect 3461 147 3477 181
rect 4245 147 4261 181
rect 4319 147 4335 181
rect 5103 147 5119 181
rect 5177 147 5193 181
rect 5961 147 5977 181
rect 6035 147 6051 181
rect 6819 147 6835 181
rect 6893 147 6909 181
rect 7677 147 7693 181
rect 7751 147 7767 181
rect 8535 147 8551 181
rect 8609 147 8625 181
rect 9393 147 9409 181
rect 9467 147 9483 181
rect 10251 147 10267 181
rect 10325 147 10341 181
rect 11109 147 11125 181
rect -11171 88 -11137 104
rect -11171 -104 -11137 -88
rect -10313 88 -10279 104
rect -10313 -104 -10279 -88
rect -9455 88 -9421 104
rect -9455 -104 -9421 -88
rect -8597 88 -8563 104
rect -8597 -104 -8563 -88
rect -7739 88 -7705 104
rect -7739 -104 -7705 -88
rect -6881 88 -6847 104
rect -6881 -104 -6847 -88
rect -6023 88 -5989 104
rect -6023 -104 -5989 -88
rect -5165 88 -5131 104
rect -5165 -104 -5131 -88
rect -4307 88 -4273 104
rect -4307 -104 -4273 -88
rect -3449 88 -3415 104
rect -3449 -104 -3415 -88
rect -2591 88 -2557 104
rect -2591 -104 -2557 -88
rect -1733 88 -1699 104
rect -1733 -104 -1699 -88
rect -875 88 -841 104
rect -875 -104 -841 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 841 88 875 104
rect 841 -104 875 -88
rect 1699 88 1733 104
rect 1699 -104 1733 -88
rect 2557 88 2591 104
rect 2557 -104 2591 -88
rect 3415 88 3449 104
rect 3415 -104 3449 -88
rect 4273 88 4307 104
rect 4273 -104 4307 -88
rect 5131 88 5165 104
rect 5131 -104 5165 -88
rect 5989 88 6023 104
rect 5989 -104 6023 -88
rect 6847 88 6881 104
rect 6847 -104 6881 -88
rect 7705 88 7739 104
rect 7705 -104 7739 -88
rect 8563 88 8597 104
rect 8563 -104 8597 -88
rect 9421 88 9455 104
rect 9421 -104 9455 -88
rect 10279 88 10313 104
rect 10279 -104 10313 -88
rect 11137 88 11171 104
rect 11137 -104 11171 -88
rect -11125 -181 -11109 -147
rect -10341 -181 -10325 -147
rect -10267 -181 -10251 -147
rect -9483 -181 -9467 -147
rect -9409 -181 -9393 -147
rect -8625 -181 -8609 -147
rect -8551 -181 -8535 -147
rect -7767 -181 -7751 -147
rect -7693 -181 -7677 -147
rect -6909 -181 -6893 -147
rect -6835 -181 -6819 -147
rect -6051 -181 -6035 -147
rect -5977 -181 -5961 -147
rect -5193 -181 -5177 -147
rect -5119 -181 -5103 -147
rect -4335 -181 -4319 -147
rect -4261 -181 -4245 -147
rect -3477 -181 -3461 -147
rect -3403 -181 -3387 -147
rect -2619 -181 -2603 -147
rect -2545 -181 -2529 -147
rect -1761 -181 -1745 -147
rect -1687 -181 -1671 -147
rect -903 -181 -887 -147
rect -829 -181 -813 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 813 -181 829 -147
rect 887 -181 903 -147
rect 1671 -181 1687 -147
rect 1745 -181 1761 -147
rect 2529 -181 2545 -147
rect 2603 -181 2619 -147
rect 3387 -181 3403 -147
rect 3461 -181 3477 -147
rect 4245 -181 4261 -147
rect 4319 -181 4335 -147
rect 5103 -181 5119 -147
rect 5177 -181 5193 -147
rect 5961 -181 5977 -147
rect 6035 -181 6051 -147
rect 6819 -181 6835 -147
rect 6893 -181 6909 -147
rect 7677 -181 7693 -147
rect 7751 -181 7767 -147
rect 8535 -181 8551 -147
rect 8609 -181 8625 -147
rect 9393 -181 9409 -147
rect 9467 -181 9483 -147
rect 10251 -181 10267 -147
rect 10325 -181 10341 -147
rect 11109 -181 11125 -147
rect -11285 -249 -11251 -187
rect 11251 -249 11285 -187
rect -11285 -283 -11189 -249
rect 11189 -283 11285 -249
<< viali >>
rect -11109 147 -10341 181
rect -10251 147 -9483 181
rect -9393 147 -8625 181
rect -8535 147 -7767 181
rect -7677 147 -6909 181
rect -6819 147 -6051 181
rect -5961 147 -5193 181
rect -5103 147 -4335 181
rect -4245 147 -3477 181
rect -3387 147 -2619 181
rect -2529 147 -1761 181
rect -1671 147 -903 181
rect -813 147 -45 181
rect 45 147 813 181
rect 903 147 1671 181
rect 1761 147 2529 181
rect 2619 147 3387 181
rect 3477 147 4245 181
rect 4335 147 5103 181
rect 5193 147 5961 181
rect 6051 147 6819 181
rect 6909 147 7677 181
rect 7767 147 8535 181
rect 8625 147 9393 181
rect 9483 147 10251 181
rect 10341 147 11109 181
rect -11171 -88 -11137 88
rect -10313 -88 -10279 88
rect -9455 -88 -9421 88
rect -8597 -88 -8563 88
rect -7739 -88 -7705 88
rect -6881 -88 -6847 88
rect -6023 -88 -5989 88
rect -5165 -88 -5131 88
rect -4307 -88 -4273 88
rect -3449 -88 -3415 88
rect -2591 -88 -2557 88
rect -1733 -88 -1699 88
rect -875 -88 -841 88
rect -17 -88 17 88
rect 841 -88 875 88
rect 1699 -88 1733 88
rect 2557 -88 2591 88
rect 3415 -88 3449 88
rect 4273 -88 4307 88
rect 5131 -88 5165 88
rect 5989 -88 6023 88
rect 6847 -88 6881 88
rect 7705 -88 7739 88
rect 8563 -88 8597 88
rect 9421 -88 9455 88
rect 10279 -88 10313 88
rect 11137 -88 11171 88
rect -11109 -181 -10341 -147
rect -10251 -181 -9483 -147
rect -9393 -181 -8625 -147
rect -8535 -181 -7767 -147
rect -7677 -181 -6909 -147
rect -6819 -181 -6051 -147
rect -5961 -181 -5193 -147
rect -5103 -181 -4335 -147
rect -4245 -181 -3477 -147
rect -3387 -181 -2619 -147
rect -2529 -181 -1761 -147
rect -1671 -181 -903 -147
rect -813 -181 -45 -147
rect 45 -181 813 -147
rect 903 -181 1671 -147
rect 1761 -181 2529 -147
rect 2619 -181 3387 -147
rect 3477 -181 4245 -147
rect 4335 -181 5103 -147
rect 5193 -181 5961 -147
rect 6051 -181 6819 -147
rect 6909 -181 7677 -147
rect 7767 -181 8535 -147
rect 8625 -181 9393 -147
rect 9483 -181 10251 -147
rect 10341 -181 11109 -147
<< metal1 >>
rect -11121 181 -10329 187
rect -11121 147 -11109 181
rect -10341 147 -10329 181
rect -11121 141 -10329 147
rect -10263 181 -9471 187
rect -10263 147 -10251 181
rect -9483 147 -9471 181
rect -10263 141 -9471 147
rect -9405 181 -8613 187
rect -9405 147 -9393 181
rect -8625 147 -8613 181
rect -9405 141 -8613 147
rect -8547 181 -7755 187
rect -8547 147 -8535 181
rect -7767 147 -7755 181
rect -8547 141 -7755 147
rect -7689 181 -6897 187
rect -7689 147 -7677 181
rect -6909 147 -6897 181
rect -7689 141 -6897 147
rect -6831 181 -6039 187
rect -6831 147 -6819 181
rect -6051 147 -6039 181
rect -6831 141 -6039 147
rect -5973 181 -5181 187
rect -5973 147 -5961 181
rect -5193 147 -5181 181
rect -5973 141 -5181 147
rect -5115 181 -4323 187
rect -5115 147 -5103 181
rect -4335 147 -4323 181
rect -5115 141 -4323 147
rect -4257 181 -3465 187
rect -4257 147 -4245 181
rect -3477 147 -3465 181
rect -4257 141 -3465 147
rect -3399 181 -2607 187
rect -3399 147 -3387 181
rect -2619 147 -2607 181
rect -3399 141 -2607 147
rect -2541 181 -1749 187
rect -2541 147 -2529 181
rect -1761 147 -1749 181
rect -2541 141 -1749 147
rect -1683 181 -891 187
rect -1683 147 -1671 181
rect -903 147 -891 181
rect -1683 141 -891 147
rect -825 181 -33 187
rect -825 147 -813 181
rect -45 147 -33 181
rect -825 141 -33 147
rect 33 181 825 187
rect 33 147 45 181
rect 813 147 825 181
rect 33 141 825 147
rect 891 181 1683 187
rect 891 147 903 181
rect 1671 147 1683 181
rect 891 141 1683 147
rect 1749 181 2541 187
rect 1749 147 1761 181
rect 2529 147 2541 181
rect 1749 141 2541 147
rect 2607 181 3399 187
rect 2607 147 2619 181
rect 3387 147 3399 181
rect 2607 141 3399 147
rect 3465 181 4257 187
rect 3465 147 3477 181
rect 4245 147 4257 181
rect 3465 141 4257 147
rect 4323 181 5115 187
rect 4323 147 4335 181
rect 5103 147 5115 181
rect 4323 141 5115 147
rect 5181 181 5973 187
rect 5181 147 5193 181
rect 5961 147 5973 181
rect 5181 141 5973 147
rect 6039 181 6831 187
rect 6039 147 6051 181
rect 6819 147 6831 181
rect 6039 141 6831 147
rect 6897 181 7689 187
rect 6897 147 6909 181
rect 7677 147 7689 181
rect 6897 141 7689 147
rect 7755 181 8547 187
rect 7755 147 7767 181
rect 8535 147 8547 181
rect 7755 141 8547 147
rect 8613 181 9405 187
rect 8613 147 8625 181
rect 9393 147 9405 181
rect 8613 141 9405 147
rect 9471 181 10263 187
rect 9471 147 9483 181
rect 10251 147 10263 181
rect 9471 141 10263 147
rect 10329 181 11121 187
rect 10329 147 10341 181
rect 11109 147 11121 181
rect 10329 141 11121 147
rect -11177 88 -11131 100
rect -11177 -88 -11171 88
rect -11137 -88 -11131 88
rect -11177 -100 -11131 -88
rect -10319 88 -10273 100
rect -10319 -88 -10313 88
rect -10279 -88 -10273 88
rect -10319 -100 -10273 -88
rect -9461 88 -9415 100
rect -9461 -88 -9455 88
rect -9421 -88 -9415 88
rect -9461 -100 -9415 -88
rect -8603 88 -8557 100
rect -8603 -88 -8597 88
rect -8563 -88 -8557 88
rect -8603 -100 -8557 -88
rect -7745 88 -7699 100
rect -7745 -88 -7739 88
rect -7705 -88 -7699 88
rect -7745 -100 -7699 -88
rect -6887 88 -6841 100
rect -6887 -88 -6881 88
rect -6847 -88 -6841 88
rect -6887 -100 -6841 -88
rect -6029 88 -5983 100
rect -6029 -88 -6023 88
rect -5989 -88 -5983 88
rect -6029 -100 -5983 -88
rect -5171 88 -5125 100
rect -5171 -88 -5165 88
rect -5131 -88 -5125 88
rect -5171 -100 -5125 -88
rect -4313 88 -4267 100
rect -4313 -88 -4307 88
rect -4273 -88 -4267 88
rect -4313 -100 -4267 -88
rect -3455 88 -3409 100
rect -3455 -88 -3449 88
rect -3415 -88 -3409 88
rect -3455 -100 -3409 -88
rect -2597 88 -2551 100
rect -2597 -88 -2591 88
rect -2557 -88 -2551 88
rect -2597 -100 -2551 -88
rect -1739 88 -1693 100
rect -1739 -88 -1733 88
rect -1699 -88 -1693 88
rect -1739 -100 -1693 -88
rect -881 88 -835 100
rect -881 -88 -875 88
rect -841 -88 -835 88
rect -881 -100 -835 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 835 88 881 100
rect 835 -88 841 88
rect 875 -88 881 88
rect 835 -100 881 -88
rect 1693 88 1739 100
rect 1693 -88 1699 88
rect 1733 -88 1739 88
rect 1693 -100 1739 -88
rect 2551 88 2597 100
rect 2551 -88 2557 88
rect 2591 -88 2597 88
rect 2551 -100 2597 -88
rect 3409 88 3455 100
rect 3409 -88 3415 88
rect 3449 -88 3455 88
rect 3409 -100 3455 -88
rect 4267 88 4313 100
rect 4267 -88 4273 88
rect 4307 -88 4313 88
rect 4267 -100 4313 -88
rect 5125 88 5171 100
rect 5125 -88 5131 88
rect 5165 -88 5171 88
rect 5125 -100 5171 -88
rect 5983 88 6029 100
rect 5983 -88 5989 88
rect 6023 -88 6029 88
rect 5983 -100 6029 -88
rect 6841 88 6887 100
rect 6841 -88 6847 88
rect 6881 -88 6887 88
rect 6841 -100 6887 -88
rect 7699 88 7745 100
rect 7699 -88 7705 88
rect 7739 -88 7745 88
rect 7699 -100 7745 -88
rect 8557 88 8603 100
rect 8557 -88 8563 88
rect 8597 -88 8603 88
rect 8557 -100 8603 -88
rect 9415 88 9461 100
rect 9415 -88 9421 88
rect 9455 -88 9461 88
rect 9415 -100 9461 -88
rect 10273 88 10319 100
rect 10273 -88 10279 88
rect 10313 -88 10319 88
rect 10273 -100 10319 -88
rect 11131 88 11177 100
rect 11131 -88 11137 88
rect 11171 -88 11177 88
rect 11131 -100 11177 -88
rect -11121 -147 -10329 -141
rect -11121 -181 -11109 -147
rect -10341 -181 -10329 -147
rect -11121 -187 -10329 -181
rect -10263 -147 -9471 -141
rect -10263 -181 -10251 -147
rect -9483 -181 -9471 -147
rect -10263 -187 -9471 -181
rect -9405 -147 -8613 -141
rect -9405 -181 -9393 -147
rect -8625 -181 -8613 -147
rect -9405 -187 -8613 -181
rect -8547 -147 -7755 -141
rect -8547 -181 -8535 -147
rect -7767 -181 -7755 -147
rect -8547 -187 -7755 -181
rect -7689 -147 -6897 -141
rect -7689 -181 -7677 -147
rect -6909 -181 -6897 -147
rect -7689 -187 -6897 -181
rect -6831 -147 -6039 -141
rect -6831 -181 -6819 -147
rect -6051 -181 -6039 -147
rect -6831 -187 -6039 -181
rect -5973 -147 -5181 -141
rect -5973 -181 -5961 -147
rect -5193 -181 -5181 -147
rect -5973 -187 -5181 -181
rect -5115 -147 -4323 -141
rect -5115 -181 -5103 -147
rect -4335 -181 -4323 -147
rect -5115 -187 -4323 -181
rect -4257 -147 -3465 -141
rect -4257 -181 -4245 -147
rect -3477 -181 -3465 -147
rect -4257 -187 -3465 -181
rect -3399 -147 -2607 -141
rect -3399 -181 -3387 -147
rect -2619 -181 -2607 -147
rect -3399 -187 -2607 -181
rect -2541 -147 -1749 -141
rect -2541 -181 -2529 -147
rect -1761 -181 -1749 -147
rect -2541 -187 -1749 -181
rect -1683 -147 -891 -141
rect -1683 -181 -1671 -147
rect -903 -181 -891 -147
rect -1683 -187 -891 -181
rect -825 -147 -33 -141
rect -825 -181 -813 -147
rect -45 -181 -33 -147
rect -825 -187 -33 -181
rect 33 -147 825 -141
rect 33 -181 45 -147
rect 813 -181 825 -147
rect 33 -187 825 -181
rect 891 -147 1683 -141
rect 891 -181 903 -147
rect 1671 -181 1683 -147
rect 891 -187 1683 -181
rect 1749 -147 2541 -141
rect 1749 -181 1761 -147
rect 2529 -181 2541 -147
rect 1749 -187 2541 -181
rect 2607 -147 3399 -141
rect 2607 -181 2619 -147
rect 3387 -181 3399 -147
rect 2607 -187 3399 -181
rect 3465 -147 4257 -141
rect 3465 -181 3477 -147
rect 4245 -181 4257 -147
rect 3465 -187 4257 -181
rect 4323 -147 5115 -141
rect 4323 -181 4335 -147
rect 5103 -181 5115 -147
rect 4323 -187 5115 -181
rect 5181 -147 5973 -141
rect 5181 -181 5193 -147
rect 5961 -181 5973 -147
rect 5181 -187 5973 -181
rect 6039 -147 6831 -141
rect 6039 -181 6051 -147
rect 6819 -181 6831 -147
rect 6039 -187 6831 -181
rect 6897 -147 7689 -141
rect 6897 -181 6909 -147
rect 7677 -181 7689 -147
rect 6897 -187 7689 -181
rect 7755 -147 8547 -141
rect 7755 -181 7767 -147
rect 8535 -181 8547 -147
rect 7755 -187 8547 -181
rect 8613 -147 9405 -141
rect 8613 -181 8625 -147
rect 9393 -181 9405 -147
rect 8613 -187 9405 -181
rect 9471 -147 10263 -141
rect 9471 -181 9483 -147
rect 10251 -181 10263 -147
rect 9471 -187 10263 -181
rect 10329 -147 11121 -141
rect 10329 -181 10341 -147
rect 11109 -181 11121 -147
rect 10329 -187 11121 -181
<< properties >>
string FIXED_BBOX -11268 -266 11268 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 4 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
