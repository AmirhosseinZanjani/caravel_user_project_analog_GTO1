magic
tech sky130A
magscale 1 2
timestamp 1699568647
<< locali >>
rect 86 2632 254 2770
rect 1366 2634 1534 2768
rect 4204 2634 4360 2768
rect 5506 2632 5674 2770
rect -94 2460 -52 2470
rect -60 2416 -52 2460
rect 5796 2460 5852 2468
rect 5796 2416 5798 2460
rect 5832 2416 5852 2460
rect 5796 2410 5852 2416
rect 76 1606 244 1744
rect 1808 1644 1862 1654
rect 1808 1610 1812 1644
rect 1860 1610 1862 1644
rect 1808 1602 1862 1610
rect 2334 1644 2388 1654
rect 2334 1610 2336 1644
rect 2384 1610 2388 1644
rect 2334 1602 2388 1610
rect 2838 1644 2902 1652
rect 2838 1610 2844 1644
rect 2892 1610 2902 1644
rect 2838 1606 2902 1610
rect 3350 1648 3424 1650
rect 3350 1614 3362 1648
rect 3410 1614 3424 1648
rect 3350 1604 3424 1614
rect 3880 1648 3946 1654
rect 3880 1614 3886 1648
rect 3934 1614 3946 1648
rect 3880 1608 3946 1614
rect 5500 1610 5668 1748
rect -100 618 1288 760
rect 75 617 1286 618
rect 1623 617 2320 654
rect 2397 617 3354 658
rect 3429 617 4124 652
rect 4461 617 5834 760
rect -102 346 46 492
rect 5688 360 5836 506
rect -80 70 14 84
rect -2 22 14 70
rect 5720 70 5838 90
rect 2790 40 2942 62
rect 2790 4 2812 40
rect 2912 4 2942 40
rect 5720 22 5744 70
rect 5822 22 5838 70
rect 5720 6 5838 22
rect 2790 -16 2942 4
<< viali >>
rect -94 2416 -60 2460
rect 5798 2416 5832 2460
rect 1812 1610 1860 1644
rect 2336 1610 2384 1644
rect 2844 1610 2892 1644
rect 3362 1614 3410 1648
rect 3886 1614 3934 1648
rect -80 22 -2 70
rect 2812 4 2912 40
rect 5744 22 5822 70
<< metal1 >>
rect 584 3012 5146 3158
rect 580 2984 5146 3012
rect 580 2676 768 2984
rect 1882 2676 2048 2984
rect 334 2634 1286 2676
rect 1624 2634 2576 2676
rect 580 2628 768 2634
rect 2648 2622 2658 2728
rect 2824 2622 2834 2728
rect 2904 2634 2914 2740
rect 3080 2634 3090 2740
rect 3676 2666 3868 2984
rect 4978 2672 5140 2984
rect 3172 2634 4116 2666
rect 4462 2634 5406 2672
rect 3676 2628 3868 2634
rect -108 2410 -98 2468
rect -42 2410 -32 2468
rect 256 2410 266 2468
rect 322 2410 332 2468
rect 770 2410 780 2468
rect 836 2410 846 2468
rect 1288 2414 1298 2472
rect 1354 2414 1364 2472
rect 1538 2418 1548 2476
rect 1604 2418 1614 2476
rect 2060 2418 2070 2476
rect 2126 2418 2136 2476
rect 2568 2418 2578 2476
rect 2634 2418 2644 2476
rect 3094 2402 3104 2582
rect 3160 2402 3170 2582
rect 3608 2408 3618 2466
rect 3674 2408 3684 2466
rect 4124 2408 4134 2466
rect 4190 2408 4200 2466
rect 4388 2410 4398 2468
rect 4454 2410 4464 2468
rect 4898 2410 4908 2468
rect 4964 2410 4974 2468
rect 5412 2412 5422 2470
rect 5478 2412 5488 2470
rect 5776 2410 5786 2468
rect 5842 2410 5852 2468
rect 0 1878 10 1936
rect 66 1878 76 1936
rect 512 1876 522 1934
rect 578 1876 588 1934
rect 1026 1878 1036 1936
rect 1092 1878 1102 1936
rect 4642 1876 4652 1934
rect 4708 1876 4718 1934
rect 5150 1882 5160 1940
rect 5216 1882 5226 1940
rect 5672 1880 5682 1938
rect 5738 1880 5748 1938
rect 1798 1810 1808 1868
rect 1864 1810 1874 1868
rect 2320 1810 2330 1868
rect 2386 1810 2396 1868
rect 2834 1800 2844 1858
rect 2900 1800 2910 1858
rect 3348 1816 3358 1874
rect 3414 1816 3424 1874
rect 3870 1812 3880 1870
rect 3936 1812 3946 1870
rect 1624 1706 2052 1740
rect 2042 1688 2052 1706
rect 2160 1706 2580 1740
rect 3172 1732 4114 1742
rect 3172 1706 3612 1732
rect 2160 1688 2170 1706
rect 3602 1680 3612 1706
rect 3720 1706 4114 1732
rect 3720 1680 3730 1706
rect 1800 1604 1810 1662
rect 1866 1604 1876 1662
rect 2324 1604 2334 1662
rect 2390 1604 2400 1662
rect 2832 1604 2842 1662
rect 2898 1604 2908 1662
rect 3348 1608 3358 1666
rect 3414 1608 3424 1666
rect 3870 1608 3880 1666
rect 3936 1608 3946 1666
rect 2416 614 2426 706
rect 2550 614 2560 706
rect 3178 614 3188 706
rect 3312 614 3322 706
rect 1798 488 1808 544
rect 1872 488 1882 544
rect 2314 488 2324 544
rect 2388 488 2398 544
rect 2834 490 2844 546
rect 2908 490 2918 546
rect 3344 492 3354 548
rect 3418 492 3428 548
rect 3860 490 3870 546
rect 3934 490 3944 546
rect 248 362 258 418
rect 322 362 332 418
rect 766 362 776 418
rect 840 362 850 418
rect 1290 362 1300 418
rect 1364 362 1374 418
rect 1544 364 1554 420
rect 1618 364 1628 420
rect 2060 362 2070 418
rect 2134 362 2144 418
rect 3604 362 3614 418
rect 3678 362 3688 418
rect 4108 370 4118 426
rect 4182 370 4192 426
rect 4372 376 4382 432
rect 4446 376 4456 432
rect 4898 374 4908 430
rect 4972 374 4982 430
rect 5418 372 5428 428
rect 5492 372 5502 428
rect -10 206 0 262
rect 64 206 74 262
rect 508 206 518 262
rect 582 206 592 262
rect 1030 204 1040 260
rect 1104 204 1114 260
rect 2568 196 2578 252
rect 2642 196 2652 252
rect 3090 204 3100 260
rect 3164 204 3174 260
rect 4640 210 4650 266
rect 4714 210 4724 266
rect 5156 208 5166 264
rect 5230 208 5240 264
rect 5668 206 5678 262
rect 5742 206 5752 262
rect 75 140 1280 142
rect -100 70 1286 140
rect 1390 90 1400 142
rect 1506 90 1516 142
rect 1623 107 2318 140
rect 3429 107 4126 142
rect 4224 88 4234 142
rect 4346 88 4356 142
rect -100 22 -80 70
rect -2 22 1286 70
rect 4446 70 5838 144
rect -100 4 1286 22
rect 2794 -2 2804 50
rect 2926 -2 2936 50
rect 4446 22 5744 70
rect 5822 22 5838 70
rect 4446 4 5838 22
<< via1 >>
rect 2658 2622 2824 2728
rect 2914 2634 3080 2740
rect -98 2460 -42 2468
rect -98 2416 -94 2460
rect -94 2416 -60 2460
rect -60 2416 -42 2460
rect -98 2410 -42 2416
rect 266 2410 322 2468
rect 780 2410 836 2468
rect 1298 2414 1354 2472
rect 1548 2418 1604 2476
rect 2070 2418 2126 2476
rect 2578 2418 2634 2476
rect 3104 2402 3160 2582
rect 3618 2408 3674 2466
rect 4134 2408 4190 2466
rect 4398 2410 4454 2468
rect 4908 2410 4964 2468
rect 5422 2412 5478 2470
rect 5786 2460 5842 2468
rect 5786 2416 5798 2460
rect 5798 2416 5832 2460
rect 5832 2416 5842 2460
rect 5786 2410 5842 2416
rect 10 1878 66 1936
rect 522 1876 578 1934
rect 1036 1878 1092 1936
rect 4652 1876 4708 1934
rect 5160 1882 5216 1940
rect 5682 1880 5738 1938
rect 1808 1810 1864 1868
rect 2330 1810 2386 1868
rect 2844 1800 2900 1858
rect 3358 1816 3414 1874
rect 3880 1812 3936 1870
rect 2052 1688 2160 1740
rect 3612 1680 3720 1732
rect 1810 1644 1866 1662
rect 1810 1610 1812 1644
rect 1812 1610 1860 1644
rect 1860 1610 1866 1644
rect 1810 1604 1866 1610
rect 2334 1644 2390 1662
rect 2334 1610 2336 1644
rect 2336 1610 2384 1644
rect 2384 1610 2390 1644
rect 2334 1604 2390 1610
rect 2842 1644 2898 1662
rect 2842 1610 2844 1644
rect 2844 1610 2892 1644
rect 2892 1610 2898 1644
rect 2842 1604 2898 1610
rect 3358 1648 3414 1666
rect 3358 1614 3362 1648
rect 3362 1614 3410 1648
rect 3410 1614 3414 1648
rect 3358 1608 3414 1614
rect 3880 1648 3936 1666
rect 3880 1614 3886 1648
rect 3886 1614 3934 1648
rect 3934 1614 3936 1648
rect 3880 1608 3936 1614
rect 2426 614 2550 706
rect 3188 614 3312 706
rect 1808 488 1872 544
rect 2324 488 2388 544
rect 2844 490 2908 546
rect 3354 492 3418 548
rect 3870 490 3934 546
rect 258 362 322 418
rect 776 362 840 418
rect 1300 362 1364 418
rect 1554 364 1618 420
rect 2070 362 2134 418
rect 3614 362 3678 418
rect 4118 370 4182 426
rect 4382 376 4446 432
rect 4908 374 4972 430
rect 5428 372 5492 428
rect 0 206 64 262
rect 518 206 582 262
rect 1040 204 1104 260
rect 2578 196 2642 252
rect 3100 204 3164 260
rect 4650 210 4714 266
rect 5166 208 5230 264
rect 5678 206 5742 262
rect 1400 90 1506 142
rect 4234 88 4346 142
rect 2804 40 2926 50
rect 2804 4 2812 40
rect 2812 4 2912 40
rect 2912 4 2926 40
rect 2804 -2 2926 4
<< metal2 >>
rect 2658 2850 3154 2912
rect 2656 2792 3154 2850
rect 2656 2738 2822 2792
rect 2914 2740 3080 2750
rect 2656 2728 2824 2738
rect 2656 2622 2658 2728
rect 2914 2632 3080 2634
rect 2656 2612 2824 2622
rect 2910 2622 3080 2632
rect 2656 2562 2822 2612
rect 3110 2592 3154 2792
rect 2910 2552 3076 2562
rect 3104 2582 3160 2592
rect 2562 2492 2678 2502
rect -98 2468 -42 2478
rect -100 2410 -98 2462
rect 266 2468 322 2478
rect -42 2410 266 2462
rect 780 2468 836 2478
rect 322 2410 780 2462
rect 1298 2472 1354 2482
rect 836 2414 1298 2462
rect 836 2410 1354 2414
rect -98 2400 -42 2410
rect 266 2400 322 2410
rect 780 2400 836 2410
rect 1298 2404 1354 2410
rect 1548 2476 1604 2486
rect 1644 2472 1772 2482
rect 1604 2418 1644 2466
rect 1548 2410 1644 2418
rect 1548 2408 1604 2410
rect 2070 2476 2126 2486
rect 1772 2418 2070 2466
rect 2126 2418 2562 2466
rect 1772 2410 2562 2418
rect 2070 2408 2126 2410
rect 2562 2396 2678 2406
rect 3102 2404 3104 2460
rect 3618 2466 3674 2476
rect 3160 2408 3618 2460
rect 4134 2466 4190 2476
rect 3948 2460 4076 2464
rect 3674 2454 4134 2460
rect 3674 2408 3948 2454
rect 3160 2404 3948 2408
rect 3104 2392 3160 2402
rect 3618 2398 3674 2404
rect 1644 2362 1772 2372
rect 4076 2408 4134 2454
rect 4076 2404 4190 2408
rect 4134 2398 4190 2404
rect 4398 2468 4454 2478
rect 4908 2468 4964 2478
rect 5422 2470 5478 2480
rect 4454 2410 4908 2468
rect 4964 2412 5422 2468
rect 5786 2468 5842 2478
rect 5478 2412 5786 2468
rect 4964 2410 5786 2412
rect 4398 2400 4454 2410
rect 4908 2400 4964 2410
rect 5422 2402 5478 2410
rect 5786 2400 5842 2410
rect 3948 2344 4076 2354
rect 5160 1946 5216 1950
rect 5682 1946 5738 1948
rect 10 1936 66 1946
rect 522 1936 578 1944
rect 1036 1936 1092 1946
rect 66 1934 1036 1936
rect 66 1878 522 1934
rect 10 1868 66 1878
rect 578 1878 1036 1934
rect 4652 1934 4708 1944
rect 5160 1940 5220 1946
rect 578 1876 580 1878
rect 522 1382 580 1876
rect 1036 1868 1092 1878
rect 1808 1868 1864 1878
rect 2330 1868 2386 1878
rect 2852 1868 2886 1900
rect 3358 1874 3414 1884
rect 1864 1810 2330 1868
rect 1808 1800 1864 1810
rect 2330 1800 2386 1810
rect 1810 1672 1862 1800
rect 2052 1740 2160 1750
rect 1810 1662 1866 1672
rect 1810 1594 1866 1604
rect 2052 1412 2160 1688
rect 2334 1672 2386 1800
rect 2844 1858 2900 1868
rect 3880 1870 3936 1880
rect 3414 1816 3880 1870
rect 3358 1812 3880 1816
rect 4708 1882 5160 1934
rect 5216 1934 5220 1940
rect 5682 1938 5742 1946
rect 5216 1882 5682 1934
rect 4708 1880 5682 1882
rect 5738 1880 5742 1938
rect 4708 1876 5742 1880
rect 4652 1866 4708 1876
rect 5160 1872 5220 1876
rect 3358 1806 3414 1812
rect 2844 1790 2900 1800
rect 2852 1672 2886 1790
rect 3360 1748 3412 1806
rect 3880 1802 3936 1812
rect 3360 1676 3414 1748
rect 3612 1740 3720 1742
rect 2334 1662 2390 1672
rect 2334 1594 2390 1604
rect 2842 1662 2898 1672
rect 2842 1594 2898 1604
rect 3358 1666 3414 1676
rect 3358 1598 3414 1608
rect 3608 1732 3720 1740
rect 3608 1680 3612 1732
rect 3608 1670 3720 1680
rect 3880 1676 3932 1802
rect 3608 1416 3716 1670
rect 3880 1666 3936 1676
rect 3880 1598 3936 1608
rect 2052 1410 2512 1412
rect 3440 1410 3716 1416
rect 1528 1382 1640 1384
rect 522 1282 1640 1382
rect 2052 1300 2578 1410
rect 1244 498 1376 508
rect 258 420 322 428
rect 776 420 840 428
rect 258 418 1244 420
rect 322 362 776 418
rect 840 362 1244 418
rect 258 352 322 362
rect 776 352 840 362
rect 1244 348 1376 358
rect 1528 420 1640 1282
rect 2410 706 2578 1300
rect 2410 614 2426 706
rect 2550 614 2578 706
rect 3178 1306 3716 1410
rect 5162 1382 5220 1872
rect 5682 1870 5742 1876
rect 3178 1304 3582 1306
rect 3178 706 3364 1304
rect 4110 1282 5224 1382
rect 4110 1252 4198 1282
rect 3178 614 3188 706
rect 3312 614 3364 706
rect 2426 604 2550 614
rect 3188 604 3312 614
rect 1808 548 3936 558
rect 1808 546 3354 548
rect 1808 544 2844 546
rect 1872 488 2324 544
rect 2388 490 2844 544
rect 2908 492 3354 546
rect 3418 546 3936 548
rect 3418 492 3870 546
rect 2908 490 3870 492
rect 3934 490 3936 546
rect 2388 488 3936 490
rect 1808 478 1872 488
rect 2324 478 2388 488
rect 2844 480 2908 488
rect 3354 482 3418 488
rect 3870 480 3934 488
rect 4112 460 4198 1252
rect 4338 498 4470 508
rect 2070 420 2134 428
rect 1528 364 1554 420
rect 1618 418 2134 420
rect 1618 364 2070 418
rect 1528 354 1640 364
rect 3614 418 3678 428
rect 2070 352 2134 362
rect 3610 362 3614 414
rect 4112 426 4194 460
rect 4112 414 4118 426
rect 3678 370 4118 414
rect 4182 370 4194 426
rect 3678 364 4194 370
rect 4908 436 4972 440
rect 5428 436 5492 438
rect 4470 430 5494 436
rect 4470 376 4908 430
rect 3678 362 4192 364
rect 3610 358 4192 362
rect 4972 428 5494 430
rect 4972 376 5428 428
rect 4908 364 4972 374
rect 5492 376 5494 428
rect 5428 362 5492 372
rect 3614 352 3678 358
rect 4338 348 4470 358
rect 0 262 64 272
rect 518 262 582 272
rect 1040 262 1104 270
rect 64 206 518 262
rect 582 260 1108 262
rect 582 206 1040 260
rect 0 196 64 206
rect 518 196 582 206
rect 1104 206 1108 260
rect 1040 194 1104 204
rect 1300 -72 1352 348
rect 2578 254 2642 262
rect 3100 260 3164 270
rect 4650 266 4714 276
rect 2578 252 3100 254
rect 2642 204 3100 252
rect 2642 196 3164 204
rect 4648 210 4650 260
rect 5166 264 5230 274
rect 4714 210 5166 260
rect 4648 208 5166 210
rect 5678 262 5742 272
rect 5230 208 5678 260
rect 4648 206 5678 208
rect 5742 206 5744 260
rect 4648 202 5744 206
rect 4650 200 4714 202
rect 5166 198 5230 202
rect 5678 196 5742 202
rect 2578 186 2642 196
rect 1400 146 1512 156
rect 1400 70 1512 80
rect 2836 60 2900 196
rect 3100 194 3164 196
rect 4234 142 4346 152
rect 4234 78 4346 88
rect 2804 50 2926 60
rect 2804 -12 2926 -2
rect 4262 -72 4318 78
rect 1300 -142 4318 -72
<< via2 >>
rect 2910 2562 3076 2622
rect 1644 2372 1772 2472
rect 2562 2476 2678 2492
rect 2562 2418 2578 2476
rect 2578 2418 2634 2476
rect 2634 2418 2678 2476
rect 2562 2406 2678 2418
rect 3948 2354 4076 2454
rect 1244 418 1376 498
rect 1244 362 1300 418
rect 1300 362 1364 418
rect 1364 362 1376 418
rect 1244 358 1376 362
rect 4338 432 4470 498
rect 4338 376 4382 432
rect 4382 376 4446 432
rect 4446 376 4470 432
rect 4338 358 4470 376
rect 1400 142 1512 146
rect 1400 90 1506 142
rect 1506 90 1512 142
rect 1400 80 1512 90
<< metal3 >>
rect 2562 2796 3082 2910
rect 2562 2497 2678 2796
rect 2908 2627 3082 2796
rect 2900 2622 3086 2627
rect 2900 2562 2910 2622
rect 3076 2562 3086 2622
rect 2900 2557 3086 2562
rect 2908 2552 3082 2557
rect 2552 2492 2688 2497
rect 1634 2472 1782 2477
rect 1634 2372 1644 2472
rect 1772 2372 1782 2472
rect 2552 2406 2562 2492
rect 2678 2406 2688 2492
rect 3944 2459 4074 2460
rect 2552 2401 2688 2406
rect 3938 2454 4086 2459
rect 1634 2367 1782 2372
rect 1644 1984 1774 2367
rect 3938 2354 3948 2454
rect 4076 2354 4086 2454
rect 3938 2349 4086 2354
rect 1264 1864 1774 1984
rect 3944 2008 4074 2349
rect 3944 1888 4460 2008
rect 1264 1252 1378 1864
rect 4342 1252 4456 1888
rect 1264 503 1376 1252
rect 4342 503 4454 1252
rect 1234 498 1386 503
rect 1234 358 1244 498
rect 1376 358 1386 498
rect 1234 353 1386 358
rect 4328 498 4480 503
rect 4328 358 4338 498
rect 4470 358 4480 498
rect 4328 353 4480 358
rect 1390 146 1522 151
rect 1390 80 1400 146
rect 1512 80 1522 146
rect 1390 75 1522 80
rect 1400 -72 1512 75
rect 4388 -72 4470 353
rect 1400 -140 4470 -72
rect 1400 -142 4460 -140
use sky130_fd_pr__nfet_01v8_ACGK3H  sky130_fd_pr__nfet_01v8_ACGK3H_0
timestamp 1699564537
transform 1 0 2868 0 1 379
box -3005 -410 3005 410
use sky130_fd_pr__pfet_01v8_564V44  sky130_fd_pr__pfet_01v8_564V44_0
timestamp 1699343385
transform 1 0 2869 0 1 2187
box -3005 -619 3005 619
<< labels >>
rlabel locali 118 2712 118 2712 1 vdd
port 2 n
rlabel metal1 1628 3074 1628 3074 1 Clk
port 1 n
rlabel metal3 1298 1256 1298 1256 1 ON
port 6 n
rlabel metal2 1528 406 1636 1384 1 NodeA1
rlabel metal2 4110 1282 5224 1382 1 NodeA2
rlabel metal3 4342 498 4454 2008 1 OP
port 5 n
rlabel locali -100 618 1288 760 1 Vss
port 0 n
rlabel locali 1623 617 2320 654 1 InP
port 3 n
rlabel locali 3429 617 4124 652 1 InN
port 4 n
<< end >>
