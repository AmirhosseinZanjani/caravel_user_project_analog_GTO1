magic
tech sky130A
magscale 1 2
timestamp 1692605656
<< error_p >>
rect -221 114 -163 120
rect -29 114 29 120
rect 163 114 221 120
rect -221 80 -209 114
rect -29 80 -17 114
rect 163 80 175 114
rect -221 74 -163 80
rect -29 74 29 80
rect 163 74 221 80
rect -317 -80 -259 -74
rect -125 -80 -67 -74
rect 67 -80 125 -74
rect 259 -80 317 -74
rect -317 -114 -305 -80
rect -125 -114 -113 -80
rect 67 -114 79 -80
rect 259 -114 271 -80
rect -317 -120 -259 -114
rect -125 -120 -67 -114
rect 67 -120 125 -114
rect 259 -120 317 -114
<< pwell >>
rect -503 -252 503 252
<< nmos >>
rect -303 -42 -273 42
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
rect 273 -42 303 42
<< ndiff >>
rect -365 30 -303 42
rect -365 -30 -353 30
rect -319 -30 -303 30
rect -365 -42 -303 -30
rect -273 30 -207 42
rect -273 -30 -257 30
rect -223 -30 -207 30
rect -273 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 273 42
rect 207 -30 223 30
rect 257 -30 273 30
rect 207 -42 273 -30
rect 303 30 365 42
rect 303 -30 319 30
rect 353 -30 365 30
rect 303 -42 365 -30
<< ndiffc >>
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
<< psubdiff >>
rect -467 182 -371 216
rect 371 182 467 216
rect -467 120 -433 182
rect 433 120 467 182
rect -467 -182 -433 -120
rect 433 -182 467 -120
rect -467 -216 -371 -182
rect 371 -216 467 -182
<< psubdiffcont >>
rect -371 182 371 216
rect -467 -120 -433 120
rect 433 -120 467 120
rect -371 -216 371 -182
<< poly >>
rect -225 114 -159 130
rect -225 80 -209 114
rect -175 80 -159 114
rect -303 42 -273 68
rect -225 64 -159 80
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -207 42 -177 64
rect -111 42 -81 68
rect -33 64 33 80
rect 159 114 225 130
rect 159 80 175 114
rect 209 80 225 114
rect -15 42 15 64
rect 81 42 111 68
rect 159 64 225 80
rect 177 42 207 64
rect 273 42 303 68
rect -303 -64 -273 -42
rect -321 -80 -255 -64
rect -207 -68 -177 -42
rect -111 -64 -81 -42
rect -321 -114 -305 -80
rect -271 -114 -255 -80
rect -321 -130 -255 -114
rect -129 -80 -63 -64
rect -15 -68 15 -42
rect 81 -64 111 -42
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect -129 -130 -63 -114
rect 63 -80 129 -64
rect 177 -68 207 -42
rect 273 -64 303 -42
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 63 -130 129 -114
rect 255 -80 321 -64
rect 255 -114 271 -80
rect 305 -114 321 -80
rect 255 -130 321 -114
<< polycont >>
rect -209 80 -175 114
rect -17 80 17 114
rect 175 80 209 114
rect -305 -114 -271 -80
rect -113 -114 -79 -80
rect 79 -114 113 -80
rect 271 -114 305 -80
<< locali >>
rect -467 182 -371 216
rect 371 182 467 216
rect -467 120 -433 182
rect 433 120 467 182
rect -225 80 -209 114
rect -175 80 -159 114
rect -33 80 -17 114
rect 17 80 33 114
rect 159 80 175 114
rect 209 80 225 114
rect -353 30 -319 46
rect -353 -46 -319 -30
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect 319 30 353 46
rect 319 -46 353 -30
rect -321 -114 -305 -80
rect -271 -114 -255 -80
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 255 -114 271 -80
rect 305 -114 321 -80
rect -467 -182 -433 -120
rect 433 -182 467 -120
rect -467 -216 -371 -182
rect 371 -216 467 -182
<< viali >>
rect -209 80 -175 114
rect -17 80 17 114
rect 175 80 209 114
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect -305 -114 -271 -80
rect -113 -114 -79 -80
rect 79 -114 113 -80
rect 271 -114 305 -80
<< metal1 >>
rect -221 114 -163 120
rect -221 80 -209 114
rect -175 80 -163 114
rect -221 74 -163 80
rect -29 114 29 120
rect -29 80 -17 114
rect 17 80 29 114
rect -29 74 29 80
rect 163 114 221 120
rect 163 80 175 114
rect 209 80 221 114
rect 163 74 221 80
rect -359 30 -313 42
rect -359 -30 -353 30
rect -319 -30 -313 30
rect -359 -42 -313 -30
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect 313 30 359 42
rect 313 -30 319 30
rect 353 -30 359 30
rect 313 -42 359 -30
rect -317 -80 -259 -74
rect -317 -114 -305 -80
rect -271 -114 -259 -80
rect -317 -120 -259 -114
rect -125 -80 -67 -74
rect -125 -114 -113 -80
rect -79 -114 -67 -80
rect -125 -120 -67 -114
rect 67 -80 125 -74
rect 67 -114 79 -80
rect 113 -114 125 -80
rect 67 -120 125 -114
rect 259 -80 317 -74
rect 259 -114 271 -80
rect 305 -114 317 -80
rect 259 -120 317 -114
<< properties >>
string FIXED_BBOX -450 -199 450 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
