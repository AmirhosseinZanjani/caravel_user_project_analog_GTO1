magic
tech sky130A
magscale 1 2
timestamp 1697806833
<< nwell >>
rect -3254 -4119 3254 4119
<< pmos >>
rect -3058 -3900 -1058 3900
rect -1000 -3900 1000 3900
rect 1058 -3900 3058 3900
<< pdiff >>
rect -3116 3888 -3058 3900
rect -3116 -3888 -3104 3888
rect -3070 -3888 -3058 3888
rect -3116 -3900 -3058 -3888
rect -1058 3888 -1000 3900
rect -1058 -3888 -1046 3888
rect -1012 -3888 -1000 3888
rect -1058 -3900 -1000 -3888
rect 1000 3888 1058 3900
rect 1000 -3888 1012 3888
rect 1046 -3888 1058 3888
rect 1000 -3900 1058 -3888
rect 3058 3888 3116 3900
rect 3058 -3888 3070 3888
rect 3104 -3888 3116 3888
rect 3058 -3900 3116 -3888
<< pdiffc >>
rect -3104 -3888 -3070 3888
rect -1046 -3888 -1012 3888
rect 1012 -3888 1046 3888
rect 3070 -3888 3104 3888
<< nsubdiff >>
rect -3218 4049 -3122 4083
rect 3122 4049 3218 4083
rect -3218 3987 -3184 4049
rect 3184 3987 3218 4049
rect -3218 -4049 -3184 -3987
rect 3184 -4049 3218 -3987
rect -3218 -4083 -3122 -4049
rect 3122 -4083 3218 -4049
<< nsubdiffcont >>
rect -3122 4049 3122 4083
rect -3218 -3987 -3184 3987
rect 3184 -3987 3218 3987
rect -3122 -4083 3122 -4049
<< poly >>
rect -3058 3981 -1058 3997
rect -3058 3947 -3042 3981
rect -1074 3947 -1058 3981
rect -3058 3900 -1058 3947
rect -1000 3981 1000 3997
rect -1000 3947 -984 3981
rect 984 3947 1000 3981
rect -1000 3900 1000 3947
rect 1058 3981 3058 3997
rect 1058 3947 1074 3981
rect 3042 3947 3058 3981
rect 1058 3900 3058 3947
rect -3058 -3947 -1058 -3900
rect -3058 -3981 -3042 -3947
rect -1074 -3981 -1058 -3947
rect -3058 -3997 -1058 -3981
rect -1000 -3947 1000 -3900
rect -1000 -3981 -984 -3947
rect 984 -3981 1000 -3947
rect -1000 -3997 1000 -3981
rect 1058 -3947 3058 -3900
rect 1058 -3981 1074 -3947
rect 3042 -3981 3058 -3947
rect 1058 -3997 3058 -3981
<< polycont >>
rect -3042 3947 -1074 3981
rect -984 3947 984 3981
rect 1074 3947 3042 3981
rect -3042 -3981 -1074 -3947
rect -984 -3981 984 -3947
rect 1074 -3981 3042 -3947
<< locali >>
rect -3218 4049 -3122 4083
rect 3122 4049 3218 4083
rect -3218 3987 -3184 4049
rect 3184 3987 3218 4049
rect -3058 3947 -3042 3981
rect -1074 3947 -1058 3981
rect -1000 3947 -984 3981
rect 984 3947 1000 3981
rect 1058 3947 1074 3981
rect 3042 3947 3058 3981
rect -3104 3888 -3070 3904
rect -3104 -3904 -3070 -3888
rect -1046 3888 -1012 3904
rect -1046 -3904 -1012 -3888
rect 1012 3888 1046 3904
rect 1012 -3904 1046 -3888
rect 3070 3888 3104 3904
rect 3070 -3904 3104 -3888
rect -3058 -3981 -3042 -3947
rect -1074 -3981 -1058 -3947
rect -1000 -3981 -984 -3947
rect 984 -3981 1000 -3947
rect 1058 -3981 1074 -3947
rect 3042 -3981 3058 -3947
rect -3218 -4049 -3184 -3987
rect 3184 -4049 3218 -3987
rect -3218 -4083 -3122 -4049
rect 3122 -4083 3218 -4049
<< viali >>
rect -3042 3947 -1074 3981
rect -984 3947 984 3981
rect 1074 3947 3042 3981
rect -3104 -3888 -3070 3888
rect -1046 -3888 -1012 3888
rect 1012 -3888 1046 3888
rect 3070 -3888 3104 3888
rect -3042 -3981 -1074 -3947
rect -984 -3981 984 -3947
rect 1074 -3981 3042 -3947
<< metal1 >>
rect -3054 3981 -1062 3987
rect -3054 3947 -3042 3981
rect -1074 3947 -1062 3981
rect -3054 3941 -1062 3947
rect -996 3981 996 3987
rect -996 3947 -984 3981
rect 984 3947 996 3981
rect -996 3941 996 3947
rect 1062 3981 3054 3987
rect 1062 3947 1074 3981
rect 3042 3947 3054 3981
rect 1062 3941 3054 3947
rect -3110 3888 -3064 3900
rect -3110 -3888 -3104 3888
rect -3070 -3888 -3064 3888
rect -3110 -3900 -3064 -3888
rect -1052 3888 -1006 3900
rect -1052 -3888 -1046 3888
rect -1012 -3888 -1006 3888
rect -1052 -3900 -1006 -3888
rect 1006 3888 1052 3900
rect 1006 -3888 1012 3888
rect 1046 -3888 1052 3888
rect 1006 -3900 1052 -3888
rect 3064 3888 3110 3900
rect 3064 -3888 3070 3888
rect 3104 -3888 3110 3888
rect 3064 -3900 3110 -3888
rect -3054 -3947 -1062 -3941
rect -3054 -3981 -3042 -3947
rect -1074 -3981 -1062 -3947
rect -3054 -3987 -1062 -3981
rect -996 -3947 996 -3941
rect -996 -3981 -984 -3947
rect 984 -3981 996 -3947
rect -996 -3987 996 -3981
rect 1062 -3947 3054 -3941
rect 1062 -3981 1074 -3947
rect 3042 -3981 3054 -3947
rect 1062 -3987 3054 -3981
<< properties >>
string FIXED_BBOX -3201 -4066 3201 4066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 39 l 10 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
