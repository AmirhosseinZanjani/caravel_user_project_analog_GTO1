magic
tech sky130A
magscale 1 2
timestamp 1681460907
<< error_p >>
rect -29 -53 29 -47
rect -29 -87 -17 -53
rect -29 -93 29 -87
<< nwell >>
rect -211 -226 211 226
<< pmos >>
rect -15 -6 15 78
<< pdiff >>
rect -73 66 -15 78
rect -73 6 -61 66
rect -27 6 -15 66
rect -73 -6 -15 6
rect 15 66 73 78
rect 15 6 27 66
rect 61 6 73 66
rect 15 -6 73 6
<< pdiffc >>
rect -61 6 -27 66
rect 27 6 61 66
<< nsubdiff >>
rect -175 156 -79 190
rect 79 156 175 190
rect -175 93 -141 156
rect 141 93 175 156
rect -175 -156 -141 -93
rect 141 -156 175 -93
rect -175 -190 -79 -156
rect 79 -190 175 -156
<< nsubdiffcont >>
rect -79 156 79 190
rect -175 -93 -141 93
rect 141 -93 175 93
rect -79 -190 79 -156
<< poly >>
rect -15 78 15 104
rect -15 -37 15 -6
rect -33 -53 33 -37
rect -33 -87 -17 -53
rect 17 -87 33 -53
rect -33 -103 33 -87
<< polycont >>
rect -17 -87 17 -53
<< locali >>
rect -175 156 -79 190
rect 79 156 175 190
rect -175 93 -141 156
rect 141 93 175 156
rect -61 66 -27 82
rect -61 -10 -27 6
rect 27 66 61 82
rect 27 -10 61 6
rect -33 -87 -17 -53
rect 17 -87 33 -53
rect -175 -156 -141 -93
rect 141 -156 175 -93
rect -175 -190 -79 -156
rect 79 -190 175 -156
<< viali >>
rect -61 6 -27 66
rect 27 6 61 66
rect -17 -87 17 -53
<< metal1 >>
rect -67 66 -21 78
rect -67 6 -61 66
rect -27 6 -21 66
rect -67 -6 -21 6
rect 21 66 67 78
rect 21 6 27 66
rect 61 6 67 66
rect 21 -6 67 6
rect -29 -53 29 -47
rect -29 -87 -17 -53
rect 17 -87 29 -53
rect -29 -93 29 -87
<< properties >>
string FIXED_BBOX -158 -173 158 173
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
