magic
tech sky130A
magscale 1 2
timestamp 1694525365
<< error_p >>
rect -671 -288 -613 -282
rect -557 -288 -499 -282
rect 499 -288 557 -282
rect 613 -288 671 -282
rect -671 -322 -659 -288
rect -557 -322 -545 -288
rect 499 -322 511 -288
rect 613 -322 625 -288
rect -671 -328 -613 -322
rect -557 -328 -499 -322
rect 499 -328 557 -322
rect 613 -328 671 -322
<< pwell >>
rect -839 -460 839 460
<< nmos >>
rect -639 -250 -609 250
rect -543 -250 -513 250
rect -447 -250 -417 250
rect -351 -250 -321 250
rect -255 -250 -225 250
rect -159 -250 -129 250
rect -63 -250 -33 250
rect 33 -250 63 250
rect 129 -250 159 250
rect 225 -250 255 250
rect 321 -250 351 250
rect 417 -250 447 250
rect 513 -250 543 250
rect 609 -250 639 250
<< ndiff >>
rect -701 238 -639 250
rect -701 -238 -689 238
rect -655 -238 -639 238
rect -701 -250 -639 -238
rect -609 238 -543 250
rect -609 -238 -593 238
rect -559 -238 -543 238
rect -609 -250 -543 -238
rect -513 238 -447 250
rect -513 -238 -497 238
rect -463 -238 -447 238
rect -513 -250 -447 -238
rect -417 238 -351 250
rect -417 -238 -401 238
rect -367 -238 -351 238
rect -417 -250 -351 -238
rect -321 238 -255 250
rect -321 -238 -305 238
rect -271 -238 -255 238
rect -321 -250 -255 -238
rect -225 238 -159 250
rect -225 -238 -209 238
rect -175 -238 -159 238
rect -225 -250 -159 -238
rect -129 238 -63 250
rect -129 -238 -113 238
rect -79 -238 -63 238
rect -129 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 129 250
rect 63 -238 79 238
rect 113 -238 129 238
rect 63 -250 129 -238
rect 159 238 225 250
rect 159 -238 175 238
rect 209 -238 225 238
rect 159 -250 225 -238
rect 255 238 321 250
rect 255 -238 271 238
rect 305 -238 321 238
rect 255 -250 321 -238
rect 351 238 417 250
rect 351 -238 367 238
rect 401 -238 417 238
rect 351 -250 417 -238
rect 447 238 513 250
rect 447 -238 463 238
rect 497 -238 513 238
rect 447 -250 513 -238
rect 543 238 609 250
rect 543 -238 559 238
rect 593 -238 609 238
rect 543 -250 609 -238
rect 639 238 701 250
rect 639 -238 655 238
rect 689 -238 701 238
rect 639 -250 701 -238
<< ndiffc >>
rect -689 -238 -655 238
rect -593 -238 -559 238
rect -497 -238 -463 238
rect -401 -238 -367 238
rect -305 -238 -271 238
rect -209 -238 -175 238
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect 175 -238 209 238
rect 271 -238 305 238
rect 367 -238 401 238
rect 463 -238 497 238
rect 559 -238 593 238
rect 655 -238 689 238
<< psubdiff >>
rect -803 390 -707 424
rect 707 390 803 424
rect -803 328 -769 390
rect 769 328 803 390
rect -803 -390 -769 -328
rect 769 -390 803 -328
rect -803 -424 -707 -390
rect 707 -424 803 -390
<< psubdiffcont >>
rect -707 390 707 424
rect -803 -328 -769 328
rect 769 -328 803 328
rect -707 -424 707 -390
<< poly >>
rect -639 250 -609 276
rect -543 250 -513 276
rect -447 250 -417 276
rect -351 250 -321 276
rect -255 250 -225 276
rect -159 250 -129 276
rect -63 250 -33 276
rect 33 250 63 276
rect 129 250 159 276
rect 225 250 255 276
rect 321 250 351 276
rect 417 250 447 276
rect 513 250 543 276
rect 609 250 639 276
rect -639 -272 -609 -250
rect -543 -272 -513 -250
rect -447 -272 -417 -250
rect -351 -272 -321 -250
rect -675 -288 -609 -272
rect -675 -322 -659 -288
rect -625 -322 -609 -288
rect -675 -338 -609 -322
rect -561 -288 -495 -272
rect -561 -322 -545 -288
rect -511 -322 -495 -288
rect -561 -338 -495 -322
rect -447 -288 -321 -272
rect -447 -322 -431 -288
rect -337 -322 -321 -288
rect -447 -338 -321 -322
rect -255 -272 -225 -250
rect -159 -272 -129 -250
rect -255 -288 -129 -272
rect -255 -322 -239 -288
rect -145 -322 -129 -288
rect -255 -338 -129 -322
rect -63 -272 -33 -250
rect 33 -272 63 -250
rect -63 -288 63 -272
rect -63 -322 -47 -288
rect 47 -322 63 -288
rect -63 -338 63 -322
rect 129 -272 159 -250
rect 225 -272 255 -250
rect 129 -288 255 -272
rect 129 -322 145 -288
rect 239 -322 255 -288
rect 129 -338 255 -322
rect 321 -272 351 -250
rect 417 -272 447 -250
rect 513 -272 543 -250
rect 609 -272 639 -250
rect 321 -288 447 -272
rect 321 -322 337 -288
rect 431 -322 447 -288
rect 321 -338 447 -322
rect 495 -288 561 -272
rect 495 -322 511 -288
rect 545 -322 561 -288
rect 495 -338 561 -322
rect 609 -288 675 -272
rect 609 -322 625 -288
rect 659 -322 675 -288
rect 609 -338 675 -322
<< polycont >>
rect -659 -322 -625 -288
rect -545 -322 -511 -288
rect -431 -322 -337 -288
rect -239 -322 -145 -288
rect -47 -322 47 -288
rect 145 -322 239 -288
rect 337 -322 431 -288
rect 511 -322 545 -288
rect 625 -322 659 -288
<< locali >>
rect -803 390 -707 424
rect 707 390 803 424
rect -803 328 -769 390
rect 769 328 803 390
rect -689 238 -655 254
rect -689 -254 -655 -238
rect -593 238 -559 254
rect -593 -254 -559 -238
rect -497 238 -463 254
rect -497 -254 -463 -238
rect -401 238 -367 254
rect -401 -254 -367 -238
rect -305 238 -271 254
rect -305 -254 -271 -238
rect -209 238 -175 254
rect -209 -254 -175 -238
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
rect 175 238 209 254
rect 175 -254 209 -238
rect 271 238 305 254
rect 271 -254 305 -238
rect 367 238 401 254
rect 367 -254 401 -238
rect 463 238 497 254
rect 463 -254 497 -238
rect 559 238 593 254
rect 559 -254 593 -238
rect 655 238 689 254
rect 655 -254 689 -238
rect -675 -322 -659 -288
rect -625 -322 -609 -288
rect -561 -322 -545 -288
rect -511 -322 -495 -288
rect -447 -322 -431 -288
rect -337 -322 -321 -288
rect -255 -322 -239 -288
rect -145 -322 -129 -288
rect -63 -322 -47 -288
rect 47 -322 63 -288
rect 129 -322 145 -288
rect 239 -322 255 -288
rect 321 -322 337 -288
rect 431 -322 447 -288
rect 495 -322 511 -288
rect 545 -322 561 -288
rect 609 -322 625 -288
rect 659 -322 675 -288
rect -803 -390 -769 -328
rect 769 -390 803 -328
rect -803 -424 -707 -390
rect 707 -424 803 -390
<< viali >>
rect -689 -238 -655 238
rect -593 -238 -559 238
rect -497 -238 -463 238
rect -401 -238 -367 238
rect -305 -238 -271 238
rect -209 -238 -175 238
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect 175 -238 209 238
rect 271 -238 305 238
rect 367 -238 401 238
rect 463 -238 497 238
rect 559 -238 593 238
rect 655 -238 689 238
rect -659 -322 -625 -288
rect -545 -322 -511 -288
rect -431 -322 -337 -288
rect -239 -322 -145 -288
rect -47 -322 47 -288
rect 145 -322 239 -288
rect 337 -322 431 -288
rect 511 -322 545 -288
rect 625 -322 659 -288
<< metal1 >>
rect -695 238 -649 250
rect -695 -238 -689 238
rect -655 -238 -649 238
rect -695 -250 -649 -238
rect -599 238 -553 250
rect -599 -238 -593 238
rect -559 -238 -553 238
rect -599 -250 -553 -238
rect -503 238 -457 250
rect -503 -238 -497 238
rect -463 -238 -457 238
rect -503 -250 -457 -238
rect -407 238 -361 250
rect -407 -238 -401 238
rect -367 -238 -361 238
rect -407 -250 -361 -238
rect -311 238 -265 250
rect -311 -238 -305 238
rect -271 -238 -265 238
rect -311 -250 -265 -238
rect -215 238 -169 250
rect -215 -238 -209 238
rect -175 -238 -169 238
rect -215 -250 -169 -238
rect -119 238 -73 250
rect -119 -238 -113 238
rect -79 -238 -73 238
rect -119 -250 -73 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 73 238 119 250
rect 73 -238 79 238
rect 113 -238 119 238
rect 73 -250 119 -238
rect 169 238 215 250
rect 169 -238 175 238
rect 209 -238 215 238
rect 169 -250 215 -238
rect 265 238 311 250
rect 265 -238 271 238
rect 305 -238 311 238
rect 265 -250 311 -238
rect 361 238 407 250
rect 361 -238 367 238
rect 401 -238 407 238
rect 361 -250 407 -238
rect 457 238 503 250
rect 457 -238 463 238
rect 497 -238 503 238
rect 457 -250 503 -238
rect 553 238 599 250
rect 553 -238 559 238
rect 593 -238 599 238
rect 553 -250 599 -238
rect 649 238 695 250
rect 649 -238 655 238
rect 689 -238 695 238
rect 649 -250 695 -238
rect -671 -288 -613 -282
rect -671 -322 -659 -288
rect -625 -322 -613 -288
rect -671 -328 -613 -322
rect -557 -288 -499 -282
rect -557 -322 -545 -288
rect -511 -322 -499 -288
rect -557 -328 -499 -322
rect -443 -288 -325 -282
rect -443 -322 -431 -288
rect -337 -322 -325 -288
rect -443 -328 -325 -322
rect -251 -288 -133 -282
rect -251 -322 -239 -288
rect -145 -322 -133 -288
rect -251 -328 -133 -322
rect -59 -288 59 -282
rect -59 -322 -47 -288
rect 47 -322 59 -288
rect -59 -328 59 -322
rect 133 -288 251 -282
rect 133 -322 145 -288
rect 239 -322 251 -288
rect 133 -328 251 -322
rect 325 -288 443 -282
rect 325 -322 337 -288
rect 431 -322 443 -288
rect 325 -328 443 -322
rect 499 -288 557 -282
rect 499 -322 511 -288
rect 545 -322 557 -288
rect 499 -328 557 -322
rect 613 -288 671 -282
rect 613 -322 625 -288
rect 659 -322 671 -288
rect 613 -328 671 -322
<< properties >>
string FIXED_BBOX -786 -407 786 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
