magic
tech sky130A
magscale 1 2
timestamp 1699543245
<< pwell >>
rect 51522 722 51574 804
<< locali >>
rect 33968 20328 68596 21104
rect 33968 20294 44066 20328
rect 44206 20294 58878 20328
rect 59018 20314 68596 20328
rect 59018 20294 68132 20314
rect 33968 20292 68132 20294
rect 33968 17748 35030 20292
rect 66662 20224 67306 20292
rect 68058 20260 68132 20292
rect 68190 20292 68596 20314
rect 68190 20260 68594 20292
rect 68058 20224 68594 20260
rect 66062 20190 68594 20224
rect 68058 19190 68594 20190
rect 68196 17748 68594 19190
rect 33968 17540 35168 17748
rect 33968 12994 35030 17540
rect 68058 16550 68594 17748
rect 68196 14360 68594 16550
rect 35980 12994 36338 13100
rect 68058 13096 68594 14360
rect 66062 13062 68594 13096
rect 66662 12994 67306 13062
rect 68058 13048 68594 13062
rect 68058 12994 68094 13048
rect 33968 12968 68094 12994
rect 68192 12968 68594 13048
rect 33968 12618 68594 12968
rect 35090 12616 68594 12618
rect 18270 5386 18528 5388
rect 84573 5386 84734 5388
rect 18270 5006 84734 5386
rect 18270 4968 43288 5006
rect 43342 4968 84734 5006
rect 18270 4967 84734 4968
rect 18270 2206 18528 4967
rect 19292 4866 19628 4967
rect 83234 4860 83522 4967
rect 84573 2974 84734 4967
rect 84452 2500 84734 2974
rect 18270 1900 18630 2206
rect 18270 690 18528 1900
rect 19304 690 19640 784
rect 31714 690 32268 794
rect 18270 658 33002 690
rect 33710 690 34264 788
rect 42108 690 42430 792
rect 44284 690 44606 792
rect 58464 690 58786 776
rect 60500 690 60822 794
rect 68704 690 69026 790
rect 33054 686 51520 690
rect 33054 658 43286 686
rect 18270 646 43286 658
rect 43344 650 51520 686
rect 51578 686 70042 690
rect 51578 652 59750 686
rect 59810 652 70042 686
rect 51578 650 70042 652
rect 70846 690 71168 790
rect 83226 690 83514 786
rect 84573 690 84734 2500
rect 70096 650 84734 690
rect 43344 646 84734 650
rect 18270 478 84734 646
<< viali >>
rect 44066 20294 44206 20328
rect 58878 20294 59018 20328
rect 68132 20260 68190 20314
rect 68094 12968 68192 13048
rect 43288 4968 43342 5006
rect 33002 658 33054 692
rect 43286 646 43344 686
rect 51520 650 51578 690
rect 59750 652 59810 686
rect 70042 650 70096 698
<< metal1 >>
rect 37988 23978 65146 24414
rect 37988 20238 38374 23978
rect 42132 22096 61014 22614
rect 42144 20246 42540 22096
rect 58816 20364 59110 20390
rect 43996 20292 44006 20364
rect 44266 20292 44276 20364
rect 58816 20292 58826 20364
rect 59086 20292 59110 20364
rect 44006 20270 44268 20292
rect 58816 20258 59110 20292
rect 37976 20224 37986 20238
rect 37254 20190 37986 20224
rect 37976 20180 37986 20190
rect 38374 20224 38384 20238
rect 42134 20226 42144 20246
rect 38374 20190 41280 20224
rect 41366 20190 42144 20226
rect 38374 20180 38384 20190
rect 42134 20188 42144 20190
rect 42532 20226 42542 20246
rect 46166 20226 46176 20248
rect 42532 20190 46176 20226
rect 46564 20226 46574 20248
rect 60618 20246 61014 22096
rect 64750 20254 65138 23978
rect 66048 20314 68206 20328
rect 66048 20260 68132 20314
rect 68190 20260 68206 20314
rect 46564 20220 51580 20226
rect 54592 20224 54602 20242
rect 46564 20190 48300 20220
rect 42532 20188 42542 20190
rect 37988 20172 38374 20180
rect 48290 20162 48300 20190
rect 48688 20190 51580 20220
rect 51656 20190 54602 20224
rect 48688 20162 48698 20190
rect 54592 20184 54602 20190
rect 54990 20224 55000 20242
rect 56724 20224 56734 20244
rect 54990 20190 56734 20224
rect 54990 20184 55000 20190
rect 56724 20186 56734 20190
rect 57122 20224 57132 20244
rect 60610 20224 60620 20246
rect 57122 20190 60620 20224
rect 57122 20186 57132 20190
rect 60610 20188 60620 20190
rect 61008 20224 61018 20246
rect 64740 20226 64750 20254
rect 61008 20190 61862 20224
rect 61946 20196 64750 20226
rect 65138 20226 65148 20254
rect 65138 20196 65976 20226
rect 61946 20190 65976 20196
rect 66048 20192 68206 20260
rect 61008 20188 61018 20190
rect 43322 16316 43332 16952
rect 43424 16316 43434 16952
rect 47436 16316 47446 16952
rect 47538 16316 47548 16952
rect 51540 16324 51550 16960
rect 51642 16324 51652 16960
rect 55674 16302 55684 16938
rect 55776 16302 55786 16938
rect 59764 16240 59774 16876
rect 59866 16240 59876 16876
rect 37174 14498 37184 15134
rect 37276 14498 37286 15134
rect 41244 14510 41254 15146
rect 41346 14510 41356 15146
rect 45388 14514 45398 15150
rect 45490 14514 45500 15150
rect 49504 14542 49514 15178
rect 49606 14542 49616 15178
rect 53620 14486 53630 15122
rect 53722 14486 53732 15122
rect 57740 14508 57750 15144
rect 57842 14508 57852 15144
rect 61852 14502 61862 15138
rect 61954 14502 61964 15138
rect 65958 14518 65968 15154
rect 66060 14518 66070 15154
rect 37170 13160 37180 13218
rect 37238 13160 37248 13218
rect 39222 13156 39232 13214
rect 39290 13156 39300 13214
rect 63914 13160 63924 13218
rect 63982 13160 63992 13218
rect 65964 13158 65974 13290
rect 66044 13158 66054 13290
rect 40374 13098 40384 13114
rect 37250 13062 40384 13098
rect 40374 13056 40384 13062
rect 40772 13098 40782 13114
rect 44280 13100 44290 13110
rect 40772 13062 41276 13098
rect 41366 13062 44290 13100
rect 40772 13056 40782 13062
rect 44280 13052 44290 13062
rect 44678 13100 44688 13110
rect 48314 13100 48324 13118
rect 44678 13062 48324 13100
rect 44678 13052 44688 13062
rect 48314 13060 48324 13062
rect 48712 13100 48722 13118
rect 48712 13062 51564 13100
rect 54600 13092 54610 13122
rect 51656 13064 54610 13092
rect 54998 13092 55008 13122
rect 58746 13092 58756 13124
rect 54998 13066 58756 13092
rect 59144 13092 59154 13124
rect 62326 13100 62336 13110
rect 59144 13066 61882 13092
rect 54998 13064 61882 13066
rect 51656 13062 61882 13064
rect 61946 13062 62336 13100
rect 48712 13060 48722 13062
rect 62326 13052 62336 13062
rect 62724 13100 62734 13110
rect 62724 13062 65984 13100
rect 62724 13052 62734 13062
rect 66100 13048 68210 13094
rect 66100 12968 68094 13048
rect 68192 12968 68210 13048
rect 66100 12960 68210 12968
rect 21208 8538 81754 9064
rect 18488 4858 20642 4992
rect 21226 4860 22236 8538
rect 25492 6284 77544 6928
rect 25492 5858 26092 6284
rect 77094 6112 77544 6284
rect 25492 5178 26086 5858
rect 25492 4860 26088 5178
rect 43276 5026 43356 5036
rect 43276 4968 43288 5026
rect 43344 4968 43356 5026
rect 43276 4956 43356 4968
rect 45419 4865 46066 4902
rect 46126 4852 46136 4916
rect 46300 4852 46308 4916
rect 50384 4864 50394 4952
rect 50650 4864 50660 4952
rect 52500 4860 52510 4948
rect 52766 4860 52776 4948
rect 56482 4848 56492 4900
rect 56592 4848 56602 4900
rect 56770 4865 57680 4898
rect 77094 4852 77546 6112
rect 77114 4850 77542 4852
rect 81090 4846 81754 8538
rect 82468 4864 84436 5002
rect 30930 4744 30940 4814
rect 31000 4744 31010 4814
rect 35048 4720 35058 4800
rect 35116 4720 35126 4800
rect 43280 4750 43290 4808
rect 43346 4750 43356 4808
rect 67974 4578 67984 4684
rect 68038 4578 68048 4684
rect 72088 4660 72098 4722
rect 72152 4660 72162 4722
rect 18590 2962 18600 3274
rect 18670 2962 18680 3274
rect 22700 2962 22710 3274
rect 22780 2962 22790 3274
rect 26796 2966 26806 3278
rect 26876 2966 26886 3278
rect 37104 3106 37114 3358
rect 37170 3106 37180 3358
rect 41220 3110 41230 3362
rect 41286 3110 41296 3362
rect 61806 3112 61816 3358
rect 61868 3112 61878 3358
rect 65906 3120 65916 3366
rect 65968 3120 65978 3366
rect 76214 2986 76224 3298
rect 76280 2986 76290 3298
rect 80324 2984 80334 3296
rect 80390 2984 80400 3296
rect 84434 2986 84444 3298
rect 84500 2986 84510 3298
rect 41190 2452 41200 2636
rect 41324 2452 41334 2636
rect 47392 2462 47402 2652
rect 47474 2462 47484 2652
rect 55608 2460 55618 2650
rect 55690 2460 55700 2650
rect 61782 2464 61792 2648
rect 61860 2464 61870 2648
rect 35050 1844 35060 2090
rect 35116 1844 35126 2090
rect 39160 1844 39170 2090
rect 39226 1844 39236 2090
rect 63852 1870 63862 2122
rect 63936 1870 63946 2122
rect 67958 1866 67968 2118
rect 68042 1866 68052 2118
rect 45336 1454 45346 1616
rect 45402 1454 45412 1616
rect 49454 1460 49464 1626
rect 49524 1460 49534 1626
rect 53578 1450 53588 1640
rect 53648 1450 53658 1640
rect 57678 1446 57688 1636
rect 57748 1446 57758 1636
rect 20610 980 20620 1148
rect 20684 980 20694 1148
rect 24752 970 24762 1138
rect 24826 970 24836 1138
rect 49452 1130 49462 1208
rect 49518 1130 49528 1208
rect 28864 962 28874 1130
rect 28938 962 28948 1130
rect 53568 1126 53578 1204
rect 53634 1126 53644 1204
rect 37102 1044 37112 1122
rect 37170 1044 37180 1122
rect 41216 1044 41226 1122
rect 41284 1044 41294 1122
rect 61804 1002 61814 1088
rect 61874 1002 61884 1088
rect 65902 1000 65912 1086
rect 65972 1000 65982 1086
rect 74144 962 74154 1076
rect 74212 962 74222 1076
rect 78262 958 78272 1072
rect 78330 958 78340 1072
rect 82370 956 82380 1070
rect 82438 956 82448 1070
rect 32990 838 33000 894
rect 33054 838 33064 894
rect 43274 856 43284 934
rect 43340 856 43350 934
rect 51510 828 51520 906
rect 51576 828 51586 906
rect 59740 840 59750 892
rect 59808 840 59818 892
rect 70030 840 70040 894
rect 70096 840 70106 894
rect 74688 805 75216 806
rect 23426 792 24020 796
rect 27760 792 28346 800
rect 18490 654 20644 788
rect 20723 755 20908 792
rect 21918 755 25150 792
rect 26286 755 28346 792
rect 28438 755 28876 792
rect 29554 774 30066 794
rect 23426 514 24020 755
rect 23420 172 24020 514
rect 27742 438 28346 755
rect 27740 176 28346 438
rect 23420 -878 24018 172
rect 27740 -688 28338 176
rect 23414 -2652 24018 -878
rect 27736 -2012 28338 -688
rect 29542 -826 30074 774
rect 35129 755 41228 792
rect 45419 755 48388 790
rect 48546 788 49452 790
rect 48546 755 49460 788
rect 53651 755 54718 790
rect 54920 755 57686 790
rect 61883 755 67972 788
rect 32976 706 33090 720
rect 32976 650 33002 706
rect 33056 650 33090 706
rect 32976 628 33090 650
rect 43276 632 43286 710
rect 43342 686 43352 710
rect 43344 646 43352 686
rect 43342 632 43352 646
rect 51482 704 51606 716
rect 70028 704 70038 708
rect 51482 690 51522 704
rect 51576 690 51606 704
rect 51482 650 51520 690
rect 51578 650 51606 690
rect 51482 640 51522 650
rect 51576 640 51606 650
rect 51482 608 51606 640
rect 59736 702 59830 704
rect 59736 650 59750 702
rect 59808 686 59830 702
rect 59810 652 59830 686
rect 59808 650 59830 652
rect 59736 628 59830 650
rect 70020 654 70038 704
rect 70094 704 70104 708
rect 70094 698 70120 704
rect 70020 650 70042 654
rect 70096 650 70120 698
rect 70020 618 70120 650
rect 72716 -316 73238 792
rect 74688 788 75222 805
rect 79084 788 79674 806
rect 74231 755 76846 788
rect 77586 755 81044 788
rect 81784 755 82372 788
rect 72712 -800 73238 -316
rect 72712 -826 73224 -800
rect 29542 -1290 73224 -826
rect 23414 -2656 24086 -2652
rect 27736 -2656 28334 -2012
rect 74688 -2292 75222 755
rect 74692 -2650 75222 -2292
rect 79084 -2650 79674 755
rect 82462 650 84430 788
rect 74692 -2654 79674 -2650
rect 74650 -2656 79674 -2654
rect 23414 -3032 79674 -2656
rect 23414 -3170 79676 -3032
rect 23414 -3174 28462 -3170
rect 74688 -3176 75222 -3170
<< via1 >>
rect 44006 20328 44266 20364
rect 44006 20294 44066 20328
rect 44066 20294 44206 20328
rect 44206 20294 44266 20328
rect 44006 20292 44266 20294
rect 58826 20328 59086 20364
rect 58826 20294 58878 20328
rect 58878 20294 59018 20328
rect 59018 20294 59086 20328
rect 58826 20292 59086 20294
rect 37986 20180 38374 20238
rect 42144 20188 42532 20246
rect 46176 20190 46564 20248
rect 48300 20162 48688 20220
rect 54602 20184 54990 20242
rect 56734 20186 57122 20244
rect 60620 20188 61008 20246
rect 64750 20196 65138 20254
rect 43332 16316 43424 16952
rect 47446 16316 47538 16952
rect 51550 16324 51642 16960
rect 55684 16302 55776 16938
rect 59774 16240 59866 16876
rect 37184 14498 37276 15134
rect 41254 14510 41346 15146
rect 45398 14514 45490 15150
rect 49514 14542 49606 15178
rect 53630 14486 53722 15122
rect 57750 14508 57842 15144
rect 61862 14502 61954 15138
rect 65968 14518 66060 15154
rect 37180 13160 37238 13218
rect 39232 13156 39290 13214
rect 63924 13160 63982 13218
rect 65974 13158 66044 13290
rect 40384 13056 40772 13114
rect 44290 13052 44678 13110
rect 48324 13060 48712 13118
rect 54610 13064 54998 13122
rect 58756 13066 59144 13124
rect 62336 13052 62724 13110
rect 43288 5006 43344 5026
rect 43288 4968 43342 5006
rect 43342 4968 43344 5006
rect 46136 4852 46300 4916
rect 50394 4864 50650 4952
rect 52510 4860 52766 4948
rect 56492 4848 56592 4900
rect 30940 4744 31000 4814
rect 35058 4720 35116 4800
rect 43290 4750 43346 4808
rect 67984 4578 68038 4684
rect 72098 4660 72152 4722
rect 18600 2962 18670 3274
rect 22710 2962 22780 3274
rect 26806 2966 26876 3278
rect 37114 3106 37170 3358
rect 41230 3110 41286 3362
rect 61816 3112 61868 3358
rect 65916 3120 65968 3366
rect 76224 2986 76280 3298
rect 80334 2984 80390 3296
rect 84444 2986 84500 3298
rect 41200 2452 41324 2636
rect 47402 2462 47474 2652
rect 55618 2460 55690 2650
rect 61792 2464 61860 2648
rect 35060 1844 35116 2090
rect 39170 1844 39226 2090
rect 63862 1870 63936 2122
rect 67968 1866 68042 2118
rect 45346 1454 45402 1616
rect 49464 1460 49524 1626
rect 53588 1450 53648 1640
rect 57688 1446 57748 1636
rect 20620 980 20684 1148
rect 24762 970 24826 1138
rect 49462 1130 49518 1208
rect 28874 962 28938 1130
rect 53578 1126 53634 1204
rect 37112 1044 37170 1122
rect 41226 1044 41284 1122
rect 61814 1002 61874 1088
rect 65912 1000 65972 1086
rect 74154 962 74212 1076
rect 78272 958 78330 1072
rect 82380 956 82438 1070
rect 33000 838 33054 894
rect 43284 856 43340 934
rect 51520 828 51576 906
rect 59750 840 59808 892
rect 70040 840 70096 894
rect 33002 692 33056 706
rect 33002 658 33054 692
rect 33054 658 33056 692
rect 33002 650 33056 658
rect 43286 686 43342 710
rect 43286 646 43342 686
rect 43286 632 43342 646
rect 51522 690 51576 704
rect 51522 650 51576 690
rect 51522 640 51576 650
rect 59750 686 59808 702
rect 59750 652 59808 686
rect 59750 650 59808 652
rect 70038 698 70094 708
rect 70038 654 70042 698
rect 70042 654 70094 698
<< metal2 >>
rect 37988 23978 65146 24414
rect 37988 20248 38374 23978
rect 42132 22096 61014 22614
rect 37986 20238 38374 20248
rect 42144 20246 42540 22096
rect 56736 21098 57112 21104
rect 46168 20716 57112 21098
rect 38374 20182 38384 20238
rect 42532 20188 42540 20246
rect 44006 20364 44266 20374
rect 37986 20170 38374 20180
rect 42144 20178 42532 20188
rect 43332 16952 43424 16962
rect 44006 16880 44266 20292
rect 46176 20258 46558 20716
rect 56736 20648 57112 20716
rect 46176 20248 46564 20258
rect 56736 20254 57116 20648
rect 58828 20374 59090 20390
rect 58826 20364 59090 20374
rect 59086 20292 59090 20364
rect 58826 20282 59090 20292
rect 54602 20242 54998 20252
rect 48300 20220 48688 20230
rect 46176 20180 46564 20190
rect 48298 20162 48300 20216
rect 54990 20184 54998 20242
rect 54602 20174 54998 20184
rect 56734 20244 57122 20254
rect 56734 20176 57122 20186
rect 48298 19702 48688 20162
rect 54604 20140 54998 20174
rect 54604 19702 54994 20140
rect 48298 19450 54994 19702
rect 47446 16952 47538 16962
rect 43424 16316 47446 16880
rect 51550 16960 51642 16970
rect 47538 16324 51550 16880
rect 55684 16938 55776 16948
rect 51642 16324 55684 16880
rect 47538 16316 55684 16324
rect 43332 16306 43424 16316
rect 47446 16306 47538 16316
rect 51550 16314 51642 16316
rect 58828 16880 59090 20282
rect 60618 20246 61014 22096
rect 60618 20188 60620 20246
rect 61008 20188 61014 20246
rect 60618 20170 61014 20188
rect 64736 20254 65146 23978
rect 64736 20196 64750 20254
rect 65138 20196 65146 20254
rect 64736 20178 65146 20196
rect 59774 16880 59866 16886
rect 55776 16876 59866 16880
rect 55776 16316 59774 16876
rect 55684 16292 55776 16302
rect 59774 16230 59866 16240
rect 49514 15178 49606 15188
rect 41254 15146 41346 15156
rect 37184 15134 37276 15144
rect 37276 14510 41254 15134
rect 45398 15150 45490 15160
rect 41346 15122 41352 15134
rect 41346 14514 45398 15122
rect 45490 14542 49514 15122
rect 65968 15154 66060 15164
rect 57750 15144 57842 15154
rect 53630 15122 53722 15132
rect 49606 14542 49692 15122
rect 45490 14514 49692 14542
rect 41346 14510 49692 14514
rect 37276 14498 49692 14510
rect 53436 14498 53630 15122
rect 37184 14488 37276 14498
rect 53722 14508 57750 15122
rect 61862 15138 61954 15148
rect 57842 14508 61862 15122
rect 53722 14502 61862 14508
rect 61954 15112 61978 15122
rect 61954 14518 65968 15112
rect 61954 14508 66060 14518
rect 61954 14502 66028 14508
rect 53722 14498 66028 14502
rect 61862 14492 61954 14498
rect 53630 14476 53722 14486
rect 48320 13936 54992 13958
rect 48320 13706 55000 13936
rect 37182 13228 37236 13250
rect 37180 13218 37238 13228
rect 37180 13150 37238 13160
rect 39232 13214 39290 13224
rect 37182 11334 37236 13150
rect 37180 9740 37240 11334
rect 39232 11254 39290 13156
rect 40384 13122 40772 13124
rect 30944 9506 31578 9508
rect 30940 9484 32000 9506
rect 30940 9258 31822 9484
rect 31996 9258 32000 9484
rect 30940 9254 32000 9258
rect 30940 4814 31000 9254
rect 31426 9252 32000 9254
rect 31822 9248 31996 9252
rect 35068 7000 35110 7004
rect 37180 7000 37244 9740
rect 39238 9502 39290 11254
rect 40382 13114 40772 13122
rect 48322 13120 48712 13706
rect 40382 13056 40384 13114
rect 40382 13046 40772 13056
rect 44290 13110 44678 13120
rect 40382 12736 40770 13046
rect 40382 11200 40772 12736
rect 44290 12646 44678 13052
rect 48324 13118 48712 13120
rect 48324 13050 48712 13060
rect 54610 13122 55000 13706
rect 65976 13300 66036 13484
rect 65974 13290 66044 13300
rect 63924 13220 63982 13228
rect 63924 13218 63986 13220
rect 63982 13160 63986 13218
rect 54998 13064 55000 13122
rect 58756 13124 59144 13134
rect 54610 13054 54998 13064
rect 58756 13056 59144 13066
rect 62336 13110 62724 13120
rect 58756 12646 59142 13056
rect 62724 13052 62736 13096
rect 62336 13042 62736 13052
rect 44288 12214 59162 12646
rect 62346 11200 62736 13042
rect 63924 11540 63986 13160
rect 65974 13148 66044 13158
rect 40382 10764 62736 11200
rect 63916 9646 63988 11540
rect 65976 10992 66036 13148
rect 39204 9488 50636 9502
rect 39298 9484 50636 9488
rect 39298 9266 50646 9484
rect 52502 9456 52752 9462
rect 63904 9456 63996 9646
rect 39204 9256 39298 9266
rect 50394 7040 50646 9266
rect 52500 9416 64000 9456
rect 52500 9194 63904 9416
rect 63998 9194 64000 9416
rect 52500 9186 64000 9194
rect 52502 7044 52752 9186
rect 63904 9184 63998 9186
rect 65974 8942 66036 10992
rect 72066 9410 72160 9420
rect 72066 9178 72160 9188
rect 35068 6792 37246 7000
rect 35068 4810 35110 6792
rect 43288 5026 43344 5036
rect 43344 4968 43346 5000
rect 43288 4958 43346 4968
rect 30940 4734 31000 4744
rect 35058 4800 35116 4810
rect 43290 4808 43346 4958
rect 50394 4952 50650 7040
rect 46136 4920 46300 4926
rect 46136 4916 46306 4920
rect 46300 4852 46306 4916
rect 52502 4958 52758 7044
rect 65974 6984 66034 8942
rect 65948 6776 68030 6984
rect 52502 4948 52766 4958
rect 52502 4944 52510 4948
rect 50394 4854 50650 4864
rect 56492 4900 56592 4910
rect 46136 4842 46306 4852
rect 52510 4850 52766 4860
rect 43290 4740 43346 4750
rect 35058 4710 35116 4720
rect 46138 4264 46306 4842
rect 56476 4848 56492 4900
rect 56592 4848 56660 4900
rect 56476 4378 56660 4848
rect 67994 4694 68028 6776
rect 72102 4732 72160 9178
rect 72098 4722 72160 4732
rect 67984 4684 68038 4694
rect 72152 4660 72158 4722
rect 72098 4654 72158 4660
rect 72098 4650 72152 4654
rect 67984 4568 68038 4578
rect 46138 4192 46308 4264
rect 56476 4192 56664 4378
rect 46138 4088 56664 4192
rect 37114 3358 37170 3368
rect 18600 3278 18670 3284
rect 22710 3278 22780 3284
rect 26806 3278 26876 3288
rect 18600 3274 26806 3278
rect 18670 2964 22710 3274
rect 18600 2952 18670 2962
rect 22780 2966 26806 3274
rect 26876 2966 26878 3278
rect 41230 3362 41286 3372
rect 37170 3110 41230 3354
rect 37170 3106 41286 3110
rect 37114 3096 37170 3106
rect 41230 3100 41286 3106
rect 61816 3358 61868 3368
rect 65916 3366 65968 3376
rect 61868 3120 65916 3358
rect 65968 3120 65970 3358
rect 61868 3112 65970 3120
rect 76224 3298 76280 3308
rect 80334 3300 80390 3306
rect 84444 3300 84500 3308
rect 61816 3102 61868 3112
rect 65916 3110 65968 3112
rect 78728 3298 84500 3300
rect 78728 3296 84444 3298
rect 76280 2986 80334 3296
rect 76224 2984 80334 2986
rect 80390 2986 84444 3296
rect 80390 2984 82004 2986
rect 76224 2982 82004 2984
rect 76224 2976 76280 2982
rect 80334 2974 80390 2982
rect 84444 2976 84500 2986
rect 22780 2964 26878 2966
rect 22710 2952 22780 2962
rect 26806 2956 26876 2964
rect 47402 2652 47474 2662
rect 55618 2652 55690 2660
rect 41200 2642 41324 2646
rect 41200 2636 47402 2642
rect 41324 2462 47402 2636
rect 47474 2650 55690 2652
rect 47474 2462 55618 2650
rect 41324 2452 49344 2462
rect 61792 2648 61860 2658
rect 55690 2464 61792 2648
rect 61860 2464 61862 2648
rect 55690 2462 61862 2464
rect 41200 2442 41324 2452
rect 55618 2450 55690 2460
rect 61792 2454 61860 2462
rect 63862 2122 63936 2132
rect 67968 2122 68042 2128
rect 35060 2092 35116 2100
rect 39170 2092 39226 2100
rect 35060 2090 39236 2092
rect 35116 1844 39170 2090
rect 39226 1844 39236 2090
rect 63936 2118 68050 2122
rect 63936 1870 67968 2118
rect 63862 1860 63936 1870
rect 68042 1870 68050 2118
rect 67968 1856 68042 1866
rect 35060 1834 35116 1844
rect 39170 1834 39226 1844
rect 45366 1648 54170 1652
rect 45366 1646 57738 1648
rect 45366 1640 57748 1646
rect 45366 1638 53588 1640
rect 45346 1626 53588 1638
rect 45346 1616 49464 1626
rect 45402 1460 49464 1616
rect 49524 1460 53588 1626
rect 45402 1458 53588 1460
rect 45346 1444 45402 1454
rect 49464 1450 49524 1458
rect 53648 1636 57748 1640
rect 53648 1458 57688 1636
rect 53588 1440 53648 1450
rect 57688 1436 57748 1446
rect 49462 1208 49518 1218
rect 53578 1208 53634 1214
rect 20620 1148 20684 1158
rect 24762 1138 24826 1148
rect 20684 980 24762 1106
rect 20620 970 20684 980
rect 28874 1130 28938 1140
rect 24826 980 28874 1106
rect 24762 960 24826 970
rect 37112 1130 37170 1132
rect 41226 1130 41284 1132
rect 49518 1204 53634 1208
rect 49518 1130 53578 1204
rect 37112 1122 41302 1130
rect 37170 1044 41226 1122
rect 41284 1044 41302 1122
rect 49462 1120 49518 1130
rect 53578 1116 53634 1126
rect 61814 1090 61874 1098
rect 65912 1090 65972 1096
rect 61814 1088 65974 1090
rect 37112 1034 37170 1044
rect 41226 1034 41284 1044
rect 61874 1086 65974 1088
rect 61874 1002 65912 1086
rect 61814 992 61874 1002
rect 65972 1002 65974 1086
rect 74154 1076 74212 1086
rect 65912 990 65972 1000
rect 28874 952 28938 962
rect 74146 962 74154 1070
rect 78272 1072 78330 1082
rect 74212 962 78272 1070
rect 74146 958 78272 962
rect 82380 1070 82438 1080
rect 78330 958 82380 1070
rect 74146 956 82380 958
rect 74146 954 82438 956
rect 74154 952 74212 954
rect 78272 948 78330 954
rect 82380 946 82438 954
rect 43284 934 43340 944
rect 33000 894 33054 904
rect 33000 828 33054 838
rect 33002 716 33054 828
rect 43284 720 43340 856
rect 51520 906 51576 916
rect 51520 818 51576 828
rect 59750 892 59808 902
rect 33002 706 33056 716
rect 43284 710 43342 720
rect 43284 652 43286 710
rect 33002 640 33056 650
rect 43286 622 43342 632
rect 51522 714 51574 818
rect 51522 704 51576 714
rect 59750 702 59808 840
rect 70040 894 70096 904
rect 70040 830 70096 840
rect 70046 718 70096 830
rect 59750 640 59808 650
rect 70038 708 70096 718
rect 70094 654 70096 708
rect 70038 644 70096 654
rect 51522 630 51576 640
<< via2 >>
rect 31822 9258 31996 9484
rect 39204 9266 39298 9488
rect 63904 9194 63998 9416
rect 72066 9188 72160 9410
<< metal3 >>
rect 31822 9492 39092 9512
rect 39194 9492 39308 9493
rect 31822 9490 39022 9492
rect 31822 9489 32008 9490
rect 31812 9484 32008 9489
rect 31812 9258 31822 9484
rect 31996 9270 32008 9484
rect 32274 9270 39022 9490
rect 39294 9488 39308 9492
rect 31996 9266 39204 9270
rect 39298 9266 39308 9488
rect 63894 9418 64008 9421
rect 31996 9258 39308 9266
rect 31812 9253 32006 9258
rect 63890 9194 63900 9418
rect 64072 9400 64082 9418
rect 72056 9410 72170 9415
rect 70072 9400 70082 9402
rect 64072 9194 70082 9400
rect 63894 9189 64008 9194
rect 70072 9184 70082 9194
rect 70418 9400 70428 9402
rect 72056 9400 72066 9410
rect 70418 9194 72066 9400
rect 70418 9184 70428 9194
rect 72056 9188 72066 9194
rect 72160 9188 72170 9410
rect 72056 9183 72170 9188
<< via3 >>
rect 32008 9270 32274 9490
rect 39022 9488 39294 9492
rect 39022 9270 39204 9488
rect 39204 9270 39294 9488
rect 63900 9416 64072 9418
rect 63900 9194 63904 9416
rect 63904 9194 63998 9416
rect 63998 9194 64072 9416
rect 70082 9184 70418 9402
<< metal4 >>
rect 24190 15490 32286 19014
rect 38894 16940 39736 16960
rect 57532 16940 67824 16950
rect 38894 16892 67824 16940
rect 38894 16266 67222 16892
rect 38894 16152 67824 16266
rect 24190 14256 32288 15490
rect 31996 9490 32288 14256
rect 31996 9270 32008 9490
rect 32274 9270 32288 9490
rect 31996 9258 32288 9270
rect 38894 9492 39736 16152
rect 57532 16144 67824 16152
rect 70098 15236 78194 19100
rect 70088 14342 78194 15236
rect 38894 9270 39022 9492
rect 39294 9270 39736 9492
rect 38894 9206 39736 9270
rect 63616 10122 64164 11036
rect 63616 9598 63808 10122
rect 64104 9598 64164 10122
rect 63616 9418 64164 9598
rect 63616 9194 63900 9418
rect 64072 9194 64164 9418
rect 70088 9403 70380 14342
rect 63616 9154 64164 9194
rect 70081 9402 70419 9403
rect 70081 9184 70082 9402
rect 70418 9184 70419 9402
rect 70081 9183 70419 9184
<< via4 >>
rect 67222 16266 68044 16892
rect 63808 9598 64104 10122
<< mimcap2 >>
rect 25102 16904 31428 18086
rect 25102 16278 30500 16904
rect 31322 16278 31428 16904
rect 25102 15164 31428 16278
rect 71010 16902 77336 18172
rect 71010 16276 71032 16902
rect 71854 16276 77336 16902
rect 71010 15250 77336 16276
<< mimcap2contact >>
rect 30500 16278 31322 16904
rect 71032 16276 71854 16902
<< metal5 >>
rect 30418 16948 64162 16958
rect 30418 16904 64166 16948
rect 30418 16278 30500 16904
rect 31322 16278 64166 16904
rect 30418 16178 64166 16278
rect 63616 10122 64166 16178
rect 67096 16902 71926 16944
rect 67096 16892 71032 16902
rect 67096 16266 67222 16892
rect 68044 16276 71032 16892
rect 71854 16276 71926 16902
rect 68044 16266 71926 16276
rect 67096 16166 71926 16266
rect 67096 16164 69738 16166
rect 63616 9598 63808 10122
rect 64104 9598 64166 10122
rect 63616 9154 64166 9598
use sky130_fd_pr__nfet_01v8_NJ4FLX  sky130_fd_pr__nfet_01v8_NJ4FLX_0
timestamp 1698072788
transform 1 0 51548 0 1 2827
box -33095 -2210 33095 2210
use sky130_fd_pr__pfet_01v8_T2K7LE  sky130_fd_pr__pfet_01v8_T2K7LE_0
timestamp 1698055914
transform 1 0 51611 0 1 16643
box -16631 -3719 16631 3719
<< labels >>
rlabel space 40382 10424 62736 11200 1 BiasP1
rlabel metal3 63998 9194 72066 9400 1 ON
rlabel metal2 65948 6776 68030 6984 1 NodeA
rlabel space 29542 -1576 73224 -826 1 BiasN2
rlabel metal2 35068 6792 37246 7000 1 NodeB
rlabel metal3 31996 9258 39092 9512 1 OP
rlabel metal1 39194 766 39194 766 1 InP
rlabel metal1 63890 766 63890 766 1 InN
rlabel metal2 37170 3106 41230 3354 1 Tail1
rlabel metal2 51544 4130 51544 4130 1 BiasTail
rlabel locali 18270 478 18270 478 3 vss
rlabel locali 33968 21102 33968 21102 1 vdd
rlabel metal2 37988 24414 37988 24414 5 BiasP1
rlabel metal2 42610 22272 42610 22272 1 BiasP2
rlabel metal1 24350 -3028 24350 -3028 1 BiasN1
rlabel metal2 44288 12214 59162 12646 1 BiasP2_uq0
rlabel metal1 32334 -1130 32334 -1130 1 BiasN2
<< end >>
