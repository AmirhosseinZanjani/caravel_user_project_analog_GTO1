magic
tech sky130A
magscale 1 2
timestamp 1697806833
<< nwell >>
rect -28979 -3719 28979 3719
<< pmos >>
rect -28783 -3500 -26783 3500
rect -26725 -3500 -24725 3500
rect -24667 -3500 -22667 3500
rect -22609 -3500 -20609 3500
rect -20551 -3500 -18551 3500
rect -18493 -3500 -16493 3500
rect -16435 -3500 -14435 3500
rect -14377 -3500 -12377 3500
rect -12319 -3500 -10319 3500
rect -10261 -3500 -8261 3500
rect -8203 -3500 -6203 3500
rect -6145 -3500 -4145 3500
rect -4087 -3500 -2087 3500
rect -2029 -3500 -29 3500
rect 29 -3500 2029 3500
rect 2087 -3500 4087 3500
rect 4145 -3500 6145 3500
rect 6203 -3500 8203 3500
rect 8261 -3500 10261 3500
rect 10319 -3500 12319 3500
rect 12377 -3500 14377 3500
rect 14435 -3500 16435 3500
rect 16493 -3500 18493 3500
rect 18551 -3500 20551 3500
rect 20609 -3500 22609 3500
rect 22667 -3500 24667 3500
rect 24725 -3500 26725 3500
rect 26783 -3500 28783 3500
<< pdiff >>
rect -28841 3488 -28783 3500
rect -28841 -3488 -28829 3488
rect -28795 -3488 -28783 3488
rect -28841 -3500 -28783 -3488
rect -26783 3488 -26725 3500
rect -26783 -3488 -26771 3488
rect -26737 -3488 -26725 3488
rect -26783 -3500 -26725 -3488
rect -24725 3488 -24667 3500
rect -24725 -3488 -24713 3488
rect -24679 -3488 -24667 3488
rect -24725 -3500 -24667 -3488
rect -22667 3488 -22609 3500
rect -22667 -3488 -22655 3488
rect -22621 -3488 -22609 3488
rect -22667 -3500 -22609 -3488
rect -20609 3488 -20551 3500
rect -20609 -3488 -20597 3488
rect -20563 -3488 -20551 3488
rect -20609 -3500 -20551 -3488
rect -18551 3488 -18493 3500
rect -18551 -3488 -18539 3488
rect -18505 -3488 -18493 3488
rect -18551 -3500 -18493 -3488
rect -16493 3488 -16435 3500
rect -16493 -3488 -16481 3488
rect -16447 -3488 -16435 3488
rect -16493 -3500 -16435 -3488
rect -14435 3488 -14377 3500
rect -14435 -3488 -14423 3488
rect -14389 -3488 -14377 3488
rect -14435 -3500 -14377 -3488
rect -12377 3488 -12319 3500
rect -12377 -3488 -12365 3488
rect -12331 -3488 -12319 3488
rect -12377 -3500 -12319 -3488
rect -10319 3488 -10261 3500
rect -10319 -3488 -10307 3488
rect -10273 -3488 -10261 3488
rect -10319 -3500 -10261 -3488
rect -8261 3488 -8203 3500
rect -8261 -3488 -8249 3488
rect -8215 -3488 -8203 3488
rect -8261 -3500 -8203 -3488
rect -6203 3488 -6145 3500
rect -6203 -3488 -6191 3488
rect -6157 -3488 -6145 3488
rect -6203 -3500 -6145 -3488
rect -4145 3488 -4087 3500
rect -4145 -3488 -4133 3488
rect -4099 -3488 -4087 3488
rect -4145 -3500 -4087 -3488
rect -2087 3488 -2029 3500
rect -2087 -3488 -2075 3488
rect -2041 -3488 -2029 3488
rect -2087 -3500 -2029 -3488
rect -29 3488 29 3500
rect -29 -3488 -17 3488
rect 17 -3488 29 3488
rect -29 -3500 29 -3488
rect 2029 3488 2087 3500
rect 2029 -3488 2041 3488
rect 2075 -3488 2087 3488
rect 2029 -3500 2087 -3488
rect 4087 3488 4145 3500
rect 4087 -3488 4099 3488
rect 4133 -3488 4145 3488
rect 4087 -3500 4145 -3488
rect 6145 3488 6203 3500
rect 6145 -3488 6157 3488
rect 6191 -3488 6203 3488
rect 6145 -3500 6203 -3488
rect 8203 3488 8261 3500
rect 8203 -3488 8215 3488
rect 8249 -3488 8261 3488
rect 8203 -3500 8261 -3488
rect 10261 3488 10319 3500
rect 10261 -3488 10273 3488
rect 10307 -3488 10319 3488
rect 10261 -3500 10319 -3488
rect 12319 3488 12377 3500
rect 12319 -3488 12331 3488
rect 12365 -3488 12377 3488
rect 12319 -3500 12377 -3488
rect 14377 3488 14435 3500
rect 14377 -3488 14389 3488
rect 14423 -3488 14435 3488
rect 14377 -3500 14435 -3488
rect 16435 3488 16493 3500
rect 16435 -3488 16447 3488
rect 16481 -3488 16493 3488
rect 16435 -3500 16493 -3488
rect 18493 3488 18551 3500
rect 18493 -3488 18505 3488
rect 18539 -3488 18551 3488
rect 18493 -3500 18551 -3488
rect 20551 3488 20609 3500
rect 20551 -3488 20563 3488
rect 20597 -3488 20609 3488
rect 20551 -3500 20609 -3488
rect 22609 3488 22667 3500
rect 22609 -3488 22621 3488
rect 22655 -3488 22667 3488
rect 22609 -3500 22667 -3488
rect 24667 3488 24725 3500
rect 24667 -3488 24679 3488
rect 24713 -3488 24725 3488
rect 24667 -3500 24725 -3488
rect 26725 3488 26783 3500
rect 26725 -3488 26737 3488
rect 26771 -3488 26783 3488
rect 26725 -3500 26783 -3488
rect 28783 3488 28841 3500
rect 28783 -3488 28795 3488
rect 28829 -3488 28841 3488
rect 28783 -3500 28841 -3488
<< pdiffc >>
rect -28829 -3488 -28795 3488
rect -26771 -3488 -26737 3488
rect -24713 -3488 -24679 3488
rect -22655 -3488 -22621 3488
rect -20597 -3488 -20563 3488
rect -18539 -3488 -18505 3488
rect -16481 -3488 -16447 3488
rect -14423 -3488 -14389 3488
rect -12365 -3488 -12331 3488
rect -10307 -3488 -10273 3488
rect -8249 -3488 -8215 3488
rect -6191 -3488 -6157 3488
rect -4133 -3488 -4099 3488
rect -2075 -3488 -2041 3488
rect -17 -3488 17 3488
rect 2041 -3488 2075 3488
rect 4099 -3488 4133 3488
rect 6157 -3488 6191 3488
rect 8215 -3488 8249 3488
rect 10273 -3488 10307 3488
rect 12331 -3488 12365 3488
rect 14389 -3488 14423 3488
rect 16447 -3488 16481 3488
rect 18505 -3488 18539 3488
rect 20563 -3488 20597 3488
rect 22621 -3488 22655 3488
rect 24679 -3488 24713 3488
rect 26737 -3488 26771 3488
rect 28795 -3488 28829 3488
<< nsubdiff >>
rect -28943 3649 -28847 3683
rect 28847 3649 28943 3683
rect -28943 3587 -28909 3649
rect 28909 3587 28943 3649
rect -28943 -3649 -28909 -3587
rect 28909 -3649 28943 -3587
rect -28943 -3683 -28847 -3649
rect 28847 -3683 28943 -3649
<< nsubdiffcont >>
rect -28847 3649 28847 3683
rect -28943 -3587 -28909 3587
rect 28909 -3587 28943 3587
rect -28847 -3683 28847 -3649
<< poly >>
rect -28783 3581 -26783 3597
rect -28783 3547 -28767 3581
rect -26799 3547 -26783 3581
rect -28783 3500 -26783 3547
rect -26725 3581 -24725 3597
rect -26725 3547 -26709 3581
rect -24741 3547 -24725 3581
rect -26725 3500 -24725 3547
rect -24667 3581 -22667 3597
rect -24667 3547 -24651 3581
rect -22683 3547 -22667 3581
rect -24667 3500 -22667 3547
rect -22609 3581 -20609 3597
rect -22609 3547 -22593 3581
rect -20625 3547 -20609 3581
rect -22609 3500 -20609 3547
rect -20551 3581 -18551 3597
rect -20551 3547 -20535 3581
rect -18567 3547 -18551 3581
rect -20551 3500 -18551 3547
rect -18493 3581 -16493 3597
rect -18493 3547 -18477 3581
rect -16509 3547 -16493 3581
rect -18493 3500 -16493 3547
rect -16435 3581 -14435 3597
rect -16435 3547 -16419 3581
rect -14451 3547 -14435 3581
rect -16435 3500 -14435 3547
rect -14377 3581 -12377 3597
rect -14377 3547 -14361 3581
rect -12393 3547 -12377 3581
rect -14377 3500 -12377 3547
rect -12319 3581 -10319 3597
rect -12319 3547 -12303 3581
rect -10335 3547 -10319 3581
rect -12319 3500 -10319 3547
rect -10261 3581 -8261 3597
rect -10261 3547 -10245 3581
rect -8277 3547 -8261 3581
rect -10261 3500 -8261 3547
rect -8203 3581 -6203 3597
rect -8203 3547 -8187 3581
rect -6219 3547 -6203 3581
rect -8203 3500 -6203 3547
rect -6145 3581 -4145 3597
rect -6145 3547 -6129 3581
rect -4161 3547 -4145 3581
rect -6145 3500 -4145 3547
rect -4087 3581 -2087 3597
rect -4087 3547 -4071 3581
rect -2103 3547 -2087 3581
rect -4087 3500 -2087 3547
rect -2029 3581 -29 3597
rect -2029 3547 -2013 3581
rect -45 3547 -29 3581
rect -2029 3500 -29 3547
rect 29 3581 2029 3597
rect 29 3547 45 3581
rect 2013 3547 2029 3581
rect 29 3500 2029 3547
rect 2087 3581 4087 3597
rect 2087 3547 2103 3581
rect 4071 3547 4087 3581
rect 2087 3500 4087 3547
rect 4145 3581 6145 3597
rect 4145 3547 4161 3581
rect 6129 3547 6145 3581
rect 4145 3500 6145 3547
rect 6203 3581 8203 3597
rect 6203 3547 6219 3581
rect 8187 3547 8203 3581
rect 6203 3500 8203 3547
rect 8261 3581 10261 3597
rect 8261 3547 8277 3581
rect 10245 3547 10261 3581
rect 8261 3500 10261 3547
rect 10319 3581 12319 3597
rect 10319 3547 10335 3581
rect 12303 3547 12319 3581
rect 10319 3500 12319 3547
rect 12377 3581 14377 3597
rect 12377 3547 12393 3581
rect 14361 3547 14377 3581
rect 12377 3500 14377 3547
rect 14435 3581 16435 3597
rect 14435 3547 14451 3581
rect 16419 3547 16435 3581
rect 14435 3500 16435 3547
rect 16493 3581 18493 3597
rect 16493 3547 16509 3581
rect 18477 3547 18493 3581
rect 16493 3500 18493 3547
rect 18551 3581 20551 3597
rect 18551 3547 18567 3581
rect 20535 3547 20551 3581
rect 18551 3500 20551 3547
rect 20609 3581 22609 3597
rect 20609 3547 20625 3581
rect 22593 3547 22609 3581
rect 20609 3500 22609 3547
rect 22667 3581 24667 3597
rect 22667 3547 22683 3581
rect 24651 3547 24667 3581
rect 22667 3500 24667 3547
rect 24725 3581 26725 3597
rect 24725 3547 24741 3581
rect 26709 3547 26725 3581
rect 24725 3500 26725 3547
rect 26783 3581 28783 3597
rect 26783 3547 26799 3581
rect 28767 3547 28783 3581
rect 26783 3500 28783 3547
rect -28783 -3547 -26783 -3500
rect -28783 -3581 -28767 -3547
rect -26799 -3581 -26783 -3547
rect -28783 -3597 -26783 -3581
rect -26725 -3547 -24725 -3500
rect -26725 -3581 -26709 -3547
rect -24741 -3581 -24725 -3547
rect -26725 -3597 -24725 -3581
rect -24667 -3547 -22667 -3500
rect -24667 -3581 -24651 -3547
rect -22683 -3581 -22667 -3547
rect -24667 -3597 -22667 -3581
rect -22609 -3547 -20609 -3500
rect -22609 -3581 -22593 -3547
rect -20625 -3581 -20609 -3547
rect -22609 -3597 -20609 -3581
rect -20551 -3547 -18551 -3500
rect -20551 -3581 -20535 -3547
rect -18567 -3581 -18551 -3547
rect -20551 -3597 -18551 -3581
rect -18493 -3547 -16493 -3500
rect -18493 -3581 -18477 -3547
rect -16509 -3581 -16493 -3547
rect -18493 -3597 -16493 -3581
rect -16435 -3547 -14435 -3500
rect -16435 -3581 -16419 -3547
rect -14451 -3581 -14435 -3547
rect -16435 -3597 -14435 -3581
rect -14377 -3547 -12377 -3500
rect -14377 -3581 -14361 -3547
rect -12393 -3581 -12377 -3547
rect -14377 -3597 -12377 -3581
rect -12319 -3547 -10319 -3500
rect -12319 -3581 -12303 -3547
rect -10335 -3581 -10319 -3547
rect -12319 -3597 -10319 -3581
rect -10261 -3547 -8261 -3500
rect -10261 -3581 -10245 -3547
rect -8277 -3581 -8261 -3547
rect -10261 -3597 -8261 -3581
rect -8203 -3547 -6203 -3500
rect -8203 -3581 -8187 -3547
rect -6219 -3581 -6203 -3547
rect -8203 -3597 -6203 -3581
rect -6145 -3547 -4145 -3500
rect -6145 -3581 -6129 -3547
rect -4161 -3581 -4145 -3547
rect -6145 -3597 -4145 -3581
rect -4087 -3547 -2087 -3500
rect -4087 -3581 -4071 -3547
rect -2103 -3581 -2087 -3547
rect -4087 -3597 -2087 -3581
rect -2029 -3547 -29 -3500
rect -2029 -3581 -2013 -3547
rect -45 -3581 -29 -3547
rect -2029 -3597 -29 -3581
rect 29 -3547 2029 -3500
rect 29 -3581 45 -3547
rect 2013 -3581 2029 -3547
rect 29 -3597 2029 -3581
rect 2087 -3547 4087 -3500
rect 2087 -3581 2103 -3547
rect 4071 -3581 4087 -3547
rect 2087 -3597 4087 -3581
rect 4145 -3547 6145 -3500
rect 4145 -3581 4161 -3547
rect 6129 -3581 6145 -3547
rect 4145 -3597 6145 -3581
rect 6203 -3547 8203 -3500
rect 6203 -3581 6219 -3547
rect 8187 -3581 8203 -3547
rect 6203 -3597 8203 -3581
rect 8261 -3547 10261 -3500
rect 8261 -3581 8277 -3547
rect 10245 -3581 10261 -3547
rect 8261 -3597 10261 -3581
rect 10319 -3547 12319 -3500
rect 10319 -3581 10335 -3547
rect 12303 -3581 12319 -3547
rect 10319 -3597 12319 -3581
rect 12377 -3547 14377 -3500
rect 12377 -3581 12393 -3547
rect 14361 -3581 14377 -3547
rect 12377 -3597 14377 -3581
rect 14435 -3547 16435 -3500
rect 14435 -3581 14451 -3547
rect 16419 -3581 16435 -3547
rect 14435 -3597 16435 -3581
rect 16493 -3547 18493 -3500
rect 16493 -3581 16509 -3547
rect 18477 -3581 18493 -3547
rect 16493 -3597 18493 -3581
rect 18551 -3547 20551 -3500
rect 18551 -3581 18567 -3547
rect 20535 -3581 20551 -3547
rect 18551 -3597 20551 -3581
rect 20609 -3547 22609 -3500
rect 20609 -3581 20625 -3547
rect 22593 -3581 22609 -3547
rect 20609 -3597 22609 -3581
rect 22667 -3547 24667 -3500
rect 22667 -3581 22683 -3547
rect 24651 -3581 24667 -3547
rect 22667 -3597 24667 -3581
rect 24725 -3547 26725 -3500
rect 24725 -3581 24741 -3547
rect 26709 -3581 26725 -3547
rect 24725 -3597 26725 -3581
rect 26783 -3547 28783 -3500
rect 26783 -3581 26799 -3547
rect 28767 -3581 28783 -3547
rect 26783 -3597 28783 -3581
<< polycont >>
rect -28767 3547 -26799 3581
rect -26709 3547 -24741 3581
rect -24651 3547 -22683 3581
rect -22593 3547 -20625 3581
rect -20535 3547 -18567 3581
rect -18477 3547 -16509 3581
rect -16419 3547 -14451 3581
rect -14361 3547 -12393 3581
rect -12303 3547 -10335 3581
rect -10245 3547 -8277 3581
rect -8187 3547 -6219 3581
rect -6129 3547 -4161 3581
rect -4071 3547 -2103 3581
rect -2013 3547 -45 3581
rect 45 3547 2013 3581
rect 2103 3547 4071 3581
rect 4161 3547 6129 3581
rect 6219 3547 8187 3581
rect 8277 3547 10245 3581
rect 10335 3547 12303 3581
rect 12393 3547 14361 3581
rect 14451 3547 16419 3581
rect 16509 3547 18477 3581
rect 18567 3547 20535 3581
rect 20625 3547 22593 3581
rect 22683 3547 24651 3581
rect 24741 3547 26709 3581
rect 26799 3547 28767 3581
rect -28767 -3581 -26799 -3547
rect -26709 -3581 -24741 -3547
rect -24651 -3581 -22683 -3547
rect -22593 -3581 -20625 -3547
rect -20535 -3581 -18567 -3547
rect -18477 -3581 -16509 -3547
rect -16419 -3581 -14451 -3547
rect -14361 -3581 -12393 -3547
rect -12303 -3581 -10335 -3547
rect -10245 -3581 -8277 -3547
rect -8187 -3581 -6219 -3547
rect -6129 -3581 -4161 -3547
rect -4071 -3581 -2103 -3547
rect -2013 -3581 -45 -3547
rect 45 -3581 2013 -3547
rect 2103 -3581 4071 -3547
rect 4161 -3581 6129 -3547
rect 6219 -3581 8187 -3547
rect 8277 -3581 10245 -3547
rect 10335 -3581 12303 -3547
rect 12393 -3581 14361 -3547
rect 14451 -3581 16419 -3547
rect 16509 -3581 18477 -3547
rect 18567 -3581 20535 -3547
rect 20625 -3581 22593 -3547
rect 22683 -3581 24651 -3547
rect 24741 -3581 26709 -3547
rect 26799 -3581 28767 -3547
<< locali >>
rect -28943 3649 -28847 3683
rect 28847 3649 28943 3683
rect -28943 3587 -28909 3649
rect 28909 3587 28943 3649
rect -28783 3547 -28767 3581
rect -26799 3547 -26783 3581
rect -26725 3547 -26709 3581
rect -24741 3547 -24725 3581
rect -24667 3547 -24651 3581
rect -22683 3547 -22667 3581
rect -22609 3547 -22593 3581
rect -20625 3547 -20609 3581
rect -20551 3547 -20535 3581
rect -18567 3547 -18551 3581
rect -18493 3547 -18477 3581
rect -16509 3547 -16493 3581
rect -16435 3547 -16419 3581
rect -14451 3547 -14435 3581
rect -14377 3547 -14361 3581
rect -12393 3547 -12377 3581
rect -12319 3547 -12303 3581
rect -10335 3547 -10319 3581
rect -10261 3547 -10245 3581
rect -8277 3547 -8261 3581
rect -8203 3547 -8187 3581
rect -6219 3547 -6203 3581
rect -6145 3547 -6129 3581
rect -4161 3547 -4145 3581
rect -4087 3547 -4071 3581
rect -2103 3547 -2087 3581
rect -2029 3547 -2013 3581
rect -45 3547 -29 3581
rect 29 3547 45 3581
rect 2013 3547 2029 3581
rect 2087 3547 2103 3581
rect 4071 3547 4087 3581
rect 4145 3547 4161 3581
rect 6129 3547 6145 3581
rect 6203 3547 6219 3581
rect 8187 3547 8203 3581
rect 8261 3547 8277 3581
rect 10245 3547 10261 3581
rect 10319 3547 10335 3581
rect 12303 3547 12319 3581
rect 12377 3547 12393 3581
rect 14361 3547 14377 3581
rect 14435 3547 14451 3581
rect 16419 3547 16435 3581
rect 16493 3547 16509 3581
rect 18477 3547 18493 3581
rect 18551 3547 18567 3581
rect 20535 3547 20551 3581
rect 20609 3547 20625 3581
rect 22593 3547 22609 3581
rect 22667 3547 22683 3581
rect 24651 3547 24667 3581
rect 24725 3547 24741 3581
rect 26709 3547 26725 3581
rect 26783 3547 26799 3581
rect 28767 3547 28783 3581
rect -28829 3488 -28795 3504
rect -28829 -3504 -28795 -3488
rect -26771 3488 -26737 3504
rect -26771 -3504 -26737 -3488
rect -24713 3488 -24679 3504
rect -24713 -3504 -24679 -3488
rect -22655 3488 -22621 3504
rect -22655 -3504 -22621 -3488
rect -20597 3488 -20563 3504
rect -20597 -3504 -20563 -3488
rect -18539 3488 -18505 3504
rect -18539 -3504 -18505 -3488
rect -16481 3488 -16447 3504
rect -16481 -3504 -16447 -3488
rect -14423 3488 -14389 3504
rect -14423 -3504 -14389 -3488
rect -12365 3488 -12331 3504
rect -12365 -3504 -12331 -3488
rect -10307 3488 -10273 3504
rect -10307 -3504 -10273 -3488
rect -8249 3488 -8215 3504
rect -8249 -3504 -8215 -3488
rect -6191 3488 -6157 3504
rect -6191 -3504 -6157 -3488
rect -4133 3488 -4099 3504
rect -4133 -3504 -4099 -3488
rect -2075 3488 -2041 3504
rect -2075 -3504 -2041 -3488
rect -17 3488 17 3504
rect -17 -3504 17 -3488
rect 2041 3488 2075 3504
rect 2041 -3504 2075 -3488
rect 4099 3488 4133 3504
rect 4099 -3504 4133 -3488
rect 6157 3488 6191 3504
rect 6157 -3504 6191 -3488
rect 8215 3488 8249 3504
rect 8215 -3504 8249 -3488
rect 10273 3488 10307 3504
rect 10273 -3504 10307 -3488
rect 12331 3488 12365 3504
rect 12331 -3504 12365 -3488
rect 14389 3488 14423 3504
rect 14389 -3504 14423 -3488
rect 16447 3488 16481 3504
rect 16447 -3504 16481 -3488
rect 18505 3488 18539 3504
rect 18505 -3504 18539 -3488
rect 20563 3488 20597 3504
rect 20563 -3504 20597 -3488
rect 22621 3488 22655 3504
rect 22621 -3504 22655 -3488
rect 24679 3488 24713 3504
rect 24679 -3504 24713 -3488
rect 26737 3488 26771 3504
rect 26737 -3504 26771 -3488
rect 28795 3488 28829 3504
rect 28795 -3504 28829 -3488
rect -28783 -3581 -28767 -3547
rect -26799 -3581 -26783 -3547
rect -26725 -3581 -26709 -3547
rect -24741 -3581 -24725 -3547
rect -24667 -3581 -24651 -3547
rect -22683 -3581 -22667 -3547
rect -22609 -3581 -22593 -3547
rect -20625 -3581 -20609 -3547
rect -20551 -3581 -20535 -3547
rect -18567 -3581 -18551 -3547
rect -18493 -3581 -18477 -3547
rect -16509 -3581 -16493 -3547
rect -16435 -3581 -16419 -3547
rect -14451 -3581 -14435 -3547
rect -14377 -3581 -14361 -3547
rect -12393 -3581 -12377 -3547
rect -12319 -3581 -12303 -3547
rect -10335 -3581 -10319 -3547
rect -10261 -3581 -10245 -3547
rect -8277 -3581 -8261 -3547
rect -8203 -3581 -8187 -3547
rect -6219 -3581 -6203 -3547
rect -6145 -3581 -6129 -3547
rect -4161 -3581 -4145 -3547
rect -4087 -3581 -4071 -3547
rect -2103 -3581 -2087 -3547
rect -2029 -3581 -2013 -3547
rect -45 -3581 -29 -3547
rect 29 -3581 45 -3547
rect 2013 -3581 2029 -3547
rect 2087 -3581 2103 -3547
rect 4071 -3581 4087 -3547
rect 4145 -3581 4161 -3547
rect 6129 -3581 6145 -3547
rect 6203 -3581 6219 -3547
rect 8187 -3581 8203 -3547
rect 8261 -3581 8277 -3547
rect 10245 -3581 10261 -3547
rect 10319 -3581 10335 -3547
rect 12303 -3581 12319 -3547
rect 12377 -3581 12393 -3547
rect 14361 -3581 14377 -3547
rect 14435 -3581 14451 -3547
rect 16419 -3581 16435 -3547
rect 16493 -3581 16509 -3547
rect 18477 -3581 18493 -3547
rect 18551 -3581 18567 -3547
rect 20535 -3581 20551 -3547
rect 20609 -3581 20625 -3547
rect 22593 -3581 22609 -3547
rect 22667 -3581 22683 -3547
rect 24651 -3581 24667 -3547
rect 24725 -3581 24741 -3547
rect 26709 -3581 26725 -3547
rect 26783 -3581 26799 -3547
rect 28767 -3581 28783 -3547
rect -28943 -3649 -28909 -3587
rect 28909 -3649 28943 -3587
rect -28943 -3683 -28847 -3649
rect 28847 -3683 28943 -3649
<< viali >>
rect -28767 3547 -26799 3581
rect -26709 3547 -24741 3581
rect -24651 3547 -22683 3581
rect -22593 3547 -20625 3581
rect -20535 3547 -18567 3581
rect -18477 3547 -16509 3581
rect -16419 3547 -14451 3581
rect -14361 3547 -12393 3581
rect -12303 3547 -10335 3581
rect -10245 3547 -8277 3581
rect -8187 3547 -6219 3581
rect -6129 3547 -4161 3581
rect -4071 3547 -2103 3581
rect -2013 3547 -45 3581
rect 45 3547 2013 3581
rect 2103 3547 4071 3581
rect 4161 3547 6129 3581
rect 6219 3547 8187 3581
rect 8277 3547 10245 3581
rect 10335 3547 12303 3581
rect 12393 3547 14361 3581
rect 14451 3547 16419 3581
rect 16509 3547 18477 3581
rect 18567 3547 20535 3581
rect 20625 3547 22593 3581
rect 22683 3547 24651 3581
rect 24741 3547 26709 3581
rect 26799 3547 28767 3581
rect -28829 -3488 -28795 3488
rect -26771 -3488 -26737 3488
rect -24713 -3488 -24679 3488
rect -22655 -3488 -22621 3488
rect -20597 -3488 -20563 3488
rect -18539 -3488 -18505 3488
rect -16481 -3488 -16447 3488
rect -14423 -3488 -14389 3488
rect -12365 -3488 -12331 3488
rect -10307 -3488 -10273 3488
rect -8249 -3488 -8215 3488
rect -6191 -3488 -6157 3488
rect -4133 -3488 -4099 3488
rect -2075 -3488 -2041 3488
rect -17 -3488 17 3488
rect 2041 -3488 2075 3488
rect 4099 -3488 4133 3488
rect 6157 -3488 6191 3488
rect 8215 -3488 8249 3488
rect 10273 -3488 10307 3488
rect 12331 -3488 12365 3488
rect 14389 -3488 14423 3488
rect 16447 -3488 16481 3488
rect 18505 -3488 18539 3488
rect 20563 -3488 20597 3488
rect 22621 -3488 22655 3488
rect 24679 -3488 24713 3488
rect 26737 -3488 26771 3488
rect 28795 -3488 28829 3488
rect -28767 -3581 -26799 -3547
rect -26709 -3581 -24741 -3547
rect -24651 -3581 -22683 -3547
rect -22593 -3581 -20625 -3547
rect -20535 -3581 -18567 -3547
rect -18477 -3581 -16509 -3547
rect -16419 -3581 -14451 -3547
rect -14361 -3581 -12393 -3547
rect -12303 -3581 -10335 -3547
rect -10245 -3581 -8277 -3547
rect -8187 -3581 -6219 -3547
rect -6129 -3581 -4161 -3547
rect -4071 -3581 -2103 -3547
rect -2013 -3581 -45 -3547
rect 45 -3581 2013 -3547
rect 2103 -3581 4071 -3547
rect 4161 -3581 6129 -3547
rect 6219 -3581 8187 -3547
rect 8277 -3581 10245 -3547
rect 10335 -3581 12303 -3547
rect 12393 -3581 14361 -3547
rect 14451 -3581 16419 -3547
rect 16509 -3581 18477 -3547
rect 18567 -3581 20535 -3547
rect 20625 -3581 22593 -3547
rect 22683 -3581 24651 -3547
rect 24741 -3581 26709 -3547
rect 26799 -3581 28767 -3547
<< metal1 >>
rect -28779 3581 -26787 3587
rect -28779 3547 -28767 3581
rect -26799 3547 -26787 3581
rect -28779 3541 -26787 3547
rect -26721 3581 -24729 3587
rect -26721 3547 -26709 3581
rect -24741 3547 -24729 3581
rect -26721 3541 -24729 3547
rect -24663 3581 -22671 3587
rect -24663 3547 -24651 3581
rect -22683 3547 -22671 3581
rect -24663 3541 -22671 3547
rect -22605 3581 -20613 3587
rect -22605 3547 -22593 3581
rect -20625 3547 -20613 3581
rect -22605 3541 -20613 3547
rect -20547 3581 -18555 3587
rect -20547 3547 -20535 3581
rect -18567 3547 -18555 3581
rect -20547 3541 -18555 3547
rect -18489 3581 -16497 3587
rect -18489 3547 -18477 3581
rect -16509 3547 -16497 3581
rect -18489 3541 -16497 3547
rect -16431 3581 -14439 3587
rect -16431 3547 -16419 3581
rect -14451 3547 -14439 3581
rect -16431 3541 -14439 3547
rect -14373 3581 -12381 3587
rect -14373 3547 -14361 3581
rect -12393 3547 -12381 3581
rect -14373 3541 -12381 3547
rect -12315 3581 -10323 3587
rect -12315 3547 -12303 3581
rect -10335 3547 -10323 3581
rect -12315 3541 -10323 3547
rect -10257 3581 -8265 3587
rect -10257 3547 -10245 3581
rect -8277 3547 -8265 3581
rect -10257 3541 -8265 3547
rect -8199 3581 -6207 3587
rect -8199 3547 -8187 3581
rect -6219 3547 -6207 3581
rect -8199 3541 -6207 3547
rect -6141 3581 -4149 3587
rect -6141 3547 -6129 3581
rect -4161 3547 -4149 3581
rect -6141 3541 -4149 3547
rect -4083 3581 -2091 3587
rect -4083 3547 -4071 3581
rect -2103 3547 -2091 3581
rect -4083 3541 -2091 3547
rect -2025 3581 -33 3587
rect -2025 3547 -2013 3581
rect -45 3547 -33 3581
rect -2025 3541 -33 3547
rect 33 3581 2025 3587
rect 33 3547 45 3581
rect 2013 3547 2025 3581
rect 33 3541 2025 3547
rect 2091 3581 4083 3587
rect 2091 3547 2103 3581
rect 4071 3547 4083 3581
rect 2091 3541 4083 3547
rect 4149 3581 6141 3587
rect 4149 3547 4161 3581
rect 6129 3547 6141 3581
rect 4149 3541 6141 3547
rect 6207 3581 8199 3587
rect 6207 3547 6219 3581
rect 8187 3547 8199 3581
rect 6207 3541 8199 3547
rect 8265 3581 10257 3587
rect 8265 3547 8277 3581
rect 10245 3547 10257 3581
rect 8265 3541 10257 3547
rect 10323 3581 12315 3587
rect 10323 3547 10335 3581
rect 12303 3547 12315 3581
rect 10323 3541 12315 3547
rect 12381 3581 14373 3587
rect 12381 3547 12393 3581
rect 14361 3547 14373 3581
rect 12381 3541 14373 3547
rect 14439 3581 16431 3587
rect 14439 3547 14451 3581
rect 16419 3547 16431 3581
rect 14439 3541 16431 3547
rect 16497 3581 18489 3587
rect 16497 3547 16509 3581
rect 18477 3547 18489 3581
rect 16497 3541 18489 3547
rect 18555 3581 20547 3587
rect 18555 3547 18567 3581
rect 20535 3547 20547 3581
rect 18555 3541 20547 3547
rect 20613 3581 22605 3587
rect 20613 3547 20625 3581
rect 22593 3547 22605 3581
rect 20613 3541 22605 3547
rect 22671 3581 24663 3587
rect 22671 3547 22683 3581
rect 24651 3547 24663 3581
rect 22671 3541 24663 3547
rect 24729 3581 26721 3587
rect 24729 3547 24741 3581
rect 26709 3547 26721 3581
rect 24729 3541 26721 3547
rect 26787 3581 28779 3587
rect 26787 3547 26799 3581
rect 28767 3547 28779 3581
rect 26787 3541 28779 3547
rect -28835 3488 -28789 3500
rect -28835 -3488 -28829 3488
rect -28795 -3488 -28789 3488
rect -28835 -3500 -28789 -3488
rect -26777 3488 -26731 3500
rect -26777 -3488 -26771 3488
rect -26737 -3488 -26731 3488
rect -26777 -3500 -26731 -3488
rect -24719 3488 -24673 3500
rect -24719 -3488 -24713 3488
rect -24679 -3488 -24673 3488
rect -24719 -3500 -24673 -3488
rect -22661 3488 -22615 3500
rect -22661 -3488 -22655 3488
rect -22621 -3488 -22615 3488
rect -22661 -3500 -22615 -3488
rect -20603 3488 -20557 3500
rect -20603 -3488 -20597 3488
rect -20563 -3488 -20557 3488
rect -20603 -3500 -20557 -3488
rect -18545 3488 -18499 3500
rect -18545 -3488 -18539 3488
rect -18505 -3488 -18499 3488
rect -18545 -3500 -18499 -3488
rect -16487 3488 -16441 3500
rect -16487 -3488 -16481 3488
rect -16447 -3488 -16441 3488
rect -16487 -3500 -16441 -3488
rect -14429 3488 -14383 3500
rect -14429 -3488 -14423 3488
rect -14389 -3488 -14383 3488
rect -14429 -3500 -14383 -3488
rect -12371 3488 -12325 3500
rect -12371 -3488 -12365 3488
rect -12331 -3488 -12325 3488
rect -12371 -3500 -12325 -3488
rect -10313 3488 -10267 3500
rect -10313 -3488 -10307 3488
rect -10273 -3488 -10267 3488
rect -10313 -3500 -10267 -3488
rect -8255 3488 -8209 3500
rect -8255 -3488 -8249 3488
rect -8215 -3488 -8209 3488
rect -8255 -3500 -8209 -3488
rect -6197 3488 -6151 3500
rect -6197 -3488 -6191 3488
rect -6157 -3488 -6151 3488
rect -6197 -3500 -6151 -3488
rect -4139 3488 -4093 3500
rect -4139 -3488 -4133 3488
rect -4099 -3488 -4093 3488
rect -4139 -3500 -4093 -3488
rect -2081 3488 -2035 3500
rect -2081 -3488 -2075 3488
rect -2041 -3488 -2035 3488
rect -2081 -3500 -2035 -3488
rect -23 3488 23 3500
rect -23 -3488 -17 3488
rect 17 -3488 23 3488
rect -23 -3500 23 -3488
rect 2035 3488 2081 3500
rect 2035 -3488 2041 3488
rect 2075 -3488 2081 3488
rect 2035 -3500 2081 -3488
rect 4093 3488 4139 3500
rect 4093 -3488 4099 3488
rect 4133 -3488 4139 3488
rect 4093 -3500 4139 -3488
rect 6151 3488 6197 3500
rect 6151 -3488 6157 3488
rect 6191 -3488 6197 3488
rect 6151 -3500 6197 -3488
rect 8209 3488 8255 3500
rect 8209 -3488 8215 3488
rect 8249 -3488 8255 3488
rect 8209 -3500 8255 -3488
rect 10267 3488 10313 3500
rect 10267 -3488 10273 3488
rect 10307 -3488 10313 3488
rect 10267 -3500 10313 -3488
rect 12325 3488 12371 3500
rect 12325 -3488 12331 3488
rect 12365 -3488 12371 3488
rect 12325 -3500 12371 -3488
rect 14383 3488 14429 3500
rect 14383 -3488 14389 3488
rect 14423 -3488 14429 3488
rect 14383 -3500 14429 -3488
rect 16441 3488 16487 3500
rect 16441 -3488 16447 3488
rect 16481 -3488 16487 3488
rect 16441 -3500 16487 -3488
rect 18499 3488 18545 3500
rect 18499 -3488 18505 3488
rect 18539 -3488 18545 3488
rect 18499 -3500 18545 -3488
rect 20557 3488 20603 3500
rect 20557 -3488 20563 3488
rect 20597 -3488 20603 3488
rect 20557 -3500 20603 -3488
rect 22615 3488 22661 3500
rect 22615 -3488 22621 3488
rect 22655 -3488 22661 3488
rect 22615 -3500 22661 -3488
rect 24673 3488 24719 3500
rect 24673 -3488 24679 3488
rect 24713 -3488 24719 3488
rect 24673 -3500 24719 -3488
rect 26731 3488 26777 3500
rect 26731 -3488 26737 3488
rect 26771 -3488 26777 3488
rect 26731 -3500 26777 -3488
rect 28789 3488 28835 3500
rect 28789 -3488 28795 3488
rect 28829 -3488 28835 3488
rect 28789 -3500 28835 -3488
rect -28779 -3547 -26787 -3541
rect -28779 -3581 -28767 -3547
rect -26799 -3581 -26787 -3547
rect -28779 -3587 -26787 -3581
rect -26721 -3547 -24729 -3541
rect -26721 -3581 -26709 -3547
rect -24741 -3581 -24729 -3547
rect -26721 -3587 -24729 -3581
rect -24663 -3547 -22671 -3541
rect -24663 -3581 -24651 -3547
rect -22683 -3581 -22671 -3547
rect -24663 -3587 -22671 -3581
rect -22605 -3547 -20613 -3541
rect -22605 -3581 -22593 -3547
rect -20625 -3581 -20613 -3547
rect -22605 -3587 -20613 -3581
rect -20547 -3547 -18555 -3541
rect -20547 -3581 -20535 -3547
rect -18567 -3581 -18555 -3547
rect -20547 -3587 -18555 -3581
rect -18489 -3547 -16497 -3541
rect -18489 -3581 -18477 -3547
rect -16509 -3581 -16497 -3547
rect -18489 -3587 -16497 -3581
rect -16431 -3547 -14439 -3541
rect -16431 -3581 -16419 -3547
rect -14451 -3581 -14439 -3547
rect -16431 -3587 -14439 -3581
rect -14373 -3547 -12381 -3541
rect -14373 -3581 -14361 -3547
rect -12393 -3581 -12381 -3547
rect -14373 -3587 -12381 -3581
rect -12315 -3547 -10323 -3541
rect -12315 -3581 -12303 -3547
rect -10335 -3581 -10323 -3547
rect -12315 -3587 -10323 -3581
rect -10257 -3547 -8265 -3541
rect -10257 -3581 -10245 -3547
rect -8277 -3581 -8265 -3547
rect -10257 -3587 -8265 -3581
rect -8199 -3547 -6207 -3541
rect -8199 -3581 -8187 -3547
rect -6219 -3581 -6207 -3547
rect -8199 -3587 -6207 -3581
rect -6141 -3547 -4149 -3541
rect -6141 -3581 -6129 -3547
rect -4161 -3581 -4149 -3547
rect -6141 -3587 -4149 -3581
rect -4083 -3547 -2091 -3541
rect -4083 -3581 -4071 -3547
rect -2103 -3581 -2091 -3547
rect -4083 -3587 -2091 -3581
rect -2025 -3547 -33 -3541
rect -2025 -3581 -2013 -3547
rect -45 -3581 -33 -3547
rect -2025 -3587 -33 -3581
rect 33 -3547 2025 -3541
rect 33 -3581 45 -3547
rect 2013 -3581 2025 -3547
rect 33 -3587 2025 -3581
rect 2091 -3547 4083 -3541
rect 2091 -3581 2103 -3547
rect 4071 -3581 4083 -3547
rect 2091 -3587 4083 -3581
rect 4149 -3547 6141 -3541
rect 4149 -3581 4161 -3547
rect 6129 -3581 6141 -3547
rect 4149 -3587 6141 -3581
rect 6207 -3547 8199 -3541
rect 6207 -3581 6219 -3547
rect 8187 -3581 8199 -3547
rect 6207 -3587 8199 -3581
rect 8265 -3547 10257 -3541
rect 8265 -3581 8277 -3547
rect 10245 -3581 10257 -3547
rect 8265 -3587 10257 -3581
rect 10323 -3547 12315 -3541
rect 10323 -3581 10335 -3547
rect 12303 -3581 12315 -3547
rect 10323 -3587 12315 -3581
rect 12381 -3547 14373 -3541
rect 12381 -3581 12393 -3547
rect 14361 -3581 14373 -3547
rect 12381 -3587 14373 -3581
rect 14439 -3547 16431 -3541
rect 14439 -3581 14451 -3547
rect 16419 -3581 16431 -3547
rect 14439 -3587 16431 -3581
rect 16497 -3547 18489 -3541
rect 16497 -3581 16509 -3547
rect 18477 -3581 18489 -3547
rect 16497 -3587 18489 -3581
rect 18555 -3547 20547 -3541
rect 18555 -3581 18567 -3547
rect 20535 -3581 20547 -3547
rect 18555 -3587 20547 -3581
rect 20613 -3547 22605 -3541
rect 20613 -3581 20625 -3547
rect 22593 -3581 22605 -3547
rect 20613 -3587 22605 -3581
rect 22671 -3547 24663 -3541
rect 22671 -3581 22683 -3547
rect 24651 -3581 24663 -3547
rect 22671 -3587 24663 -3581
rect 24729 -3547 26721 -3541
rect 24729 -3581 24741 -3547
rect 26709 -3581 26721 -3547
rect 24729 -3587 26721 -3581
rect 26787 -3547 28779 -3541
rect 26787 -3581 26799 -3547
rect 28767 -3581 28779 -3547
rect 26787 -3587 28779 -3581
<< properties >>
string FIXED_BBOX -28926 -3666 28926 3666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 35 l 10 m 1 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
