magic
tech sky130A
magscale 1 2
timestamp 1699485026
<< pwell >>
rect -33095 -2210 33095 2210
<< nmos >>
rect -32899 -2000 -30899 2000
rect -30841 -2000 -28841 2000
rect -28783 -2000 -26783 2000
rect -26725 -2000 -24725 2000
rect -24667 -2000 -22667 2000
rect -22609 -2000 -20609 2000
rect -20551 -2000 -18551 2000
rect -18493 -2000 -16493 2000
rect -16435 -2000 -14435 2000
rect -14377 -2000 -12377 2000
rect -12319 -2000 -10319 2000
rect -10261 -2000 -8261 2000
rect -8203 -2000 -6203 2000
rect -6145 -2000 -4145 2000
rect -4087 -2000 -2087 2000
rect -2029 -2000 -29 2000
rect 29 -2000 2029 2000
rect 2087 -2000 4087 2000
rect 4145 -2000 6145 2000
rect 6203 -2000 8203 2000
rect 8261 -2000 10261 2000
rect 10319 -2000 12319 2000
rect 12377 -2000 14377 2000
rect 14435 -2000 16435 2000
rect 16493 -2000 18493 2000
rect 18551 -2000 20551 2000
rect 20609 -2000 22609 2000
rect 22667 -2000 24667 2000
rect 24725 -2000 26725 2000
rect 26783 -2000 28783 2000
rect 28841 -2000 30841 2000
rect 30899 -2000 32899 2000
<< ndiff >>
rect -32957 1988 -32899 2000
rect -32957 -1988 -32945 1988
rect -32911 -1988 -32899 1988
rect -32957 -2000 -32899 -1988
rect -30899 1988 -30841 2000
rect -30899 -1988 -30887 1988
rect -30853 -1988 -30841 1988
rect -30899 -2000 -30841 -1988
rect -28841 1988 -28783 2000
rect -28841 -1988 -28829 1988
rect -28795 -1988 -28783 1988
rect -28841 -2000 -28783 -1988
rect -26783 1988 -26725 2000
rect -26783 -1988 -26771 1988
rect -26737 -1988 -26725 1988
rect -26783 -2000 -26725 -1988
rect -24725 1988 -24667 2000
rect -24725 -1988 -24713 1988
rect -24679 -1988 -24667 1988
rect -24725 -2000 -24667 -1988
rect -22667 1988 -22609 2000
rect -22667 -1988 -22655 1988
rect -22621 -1988 -22609 1988
rect -22667 -2000 -22609 -1988
rect -20609 1988 -20551 2000
rect -20609 -1988 -20597 1988
rect -20563 -1988 -20551 1988
rect -20609 -2000 -20551 -1988
rect -18551 1988 -18493 2000
rect -18551 -1988 -18539 1988
rect -18505 -1988 -18493 1988
rect -18551 -2000 -18493 -1988
rect -16493 1988 -16435 2000
rect -16493 -1988 -16481 1988
rect -16447 -1988 -16435 1988
rect -16493 -2000 -16435 -1988
rect -14435 1988 -14377 2000
rect -14435 -1988 -14423 1988
rect -14389 -1988 -14377 1988
rect -14435 -2000 -14377 -1988
rect -12377 1988 -12319 2000
rect -12377 -1988 -12365 1988
rect -12331 -1988 -12319 1988
rect -12377 -2000 -12319 -1988
rect -10319 1988 -10261 2000
rect -10319 -1988 -10307 1988
rect -10273 -1988 -10261 1988
rect -10319 -2000 -10261 -1988
rect -8261 1988 -8203 2000
rect -8261 -1988 -8249 1988
rect -8215 -1988 -8203 1988
rect -8261 -2000 -8203 -1988
rect -6203 1988 -6145 2000
rect -6203 -1988 -6191 1988
rect -6157 -1988 -6145 1988
rect -6203 -2000 -6145 -1988
rect -4145 1988 -4087 2000
rect -4145 -1988 -4133 1988
rect -4099 -1988 -4087 1988
rect -4145 -2000 -4087 -1988
rect -2087 1988 -2029 2000
rect -2087 -1988 -2075 1988
rect -2041 -1988 -2029 1988
rect -2087 -2000 -2029 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 2029 1988 2087 2000
rect 2029 -1988 2041 1988
rect 2075 -1988 2087 1988
rect 2029 -2000 2087 -1988
rect 4087 1988 4145 2000
rect 4087 -1988 4099 1988
rect 4133 -1988 4145 1988
rect 4087 -2000 4145 -1988
rect 6145 1988 6203 2000
rect 6145 -1988 6157 1988
rect 6191 -1988 6203 1988
rect 6145 -2000 6203 -1988
rect 8203 1988 8261 2000
rect 8203 -1988 8215 1988
rect 8249 -1988 8261 1988
rect 8203 -2000 8261 -1988
rect 10261 1988 10319 2000
rect 10261 -1988 10273 1988
rect 10307 -1988 10319 1988
rect 10261 -2000 10319 -1988
rect 12319 1988 12377 2000
rect 12319 -1988 12331 1988
rect 12365 -1988 12377 1988
rect 12319 -2000 12377 -1988
rect 14377 1988 14435 2000
rect 14377 -1988 14389 1988
rect 14423 -1988 14435 1988
rect 14377 -2000 14435 -1988
rect 16435 1988 16493 2000
rect 16435 -1988 16447 1988
rect 16481 -1988 16493 1988
rect 16435 -2000 16493 -1988
rect 18493 1988 18551 2000
rect 18493 -1988 18505 1988
rect 18539 -1988 18551 1988
rect 18493 -2000 18551 -1988
rect 20551 1988 20609 2000
rect 20551 -1988 20563 1988
rect 20597 -1988 20609 1988
rect 20551 -2000 20609 -1988
rect 22609 1988 22667 2000
rect 22609 -1988 22621 1988
rect 22655 -1988 22667 1988
rect 22609 -2000 22667 -1988
rect 24667 1988 24725 2000
rect 24667 -1988 24679 1988
rect 24713 -1988 24725 1988
rect 24667 -2000 24725 -1988
rect 26725 1988 26783 2000
rect 26725 -1988 26737 1988
rect 26771 -1988 26783 1988
rect 26725 -2000 26783 -1988
rect 28783 1988 28841 2000
rect 28783 -1988 28795 1988
rect 28829 -1988 28841 1988
rect 28783 -2000 28841 -1988
rect 30841 1988 30899 2000
rect 30841 -1988 30853 1988
rect 30887 -1988 30899 1988
rect 30841 -2000 30899 -1988
rect 32899 1988 32957 2000
rect 32899 -1988 32911 1988
rect 32945 -1988 32957 1988
rect 32899 -2000 32957 -1988
<< ndiffc >>
rect -32945 -1988 -32911 1988
rect -30887 -1988 -30853 1988
rect -28829 -1988 -28795 1988
rect -26771 -1988 -26737 1988
rect -24713 -1988 -24679 1988
rect -22655 -1988 -22621 1988
rect -20597 -1988 -20563 1988
rect -18539 -1988 -18505 1988
rect -16481 -1988 -16447 1988
rect -14423 -1988 -14389 1988
rect -12365 -1988 -12331 1988
rect -10307 -1988 -10273 1988
rect -8249 -1988 -8215 1988
rect -6191 -1988 -6157 1988
rect -4133 -1988 -4099 1988
rect -2075 -1988 -2041 1988
rect -17 -1988 17 1988
rect 2041 -1988 2075 1988
rect 4099 -1988 4133 1988
rect 6157 -1988 6191 1988
rect 8215 -1988 8249 1988
rect 10273 -1988 10307 1988
rect 12331 -1988 12365 1988
rect 14389 -1988 14423 1988
rect 16447 -1988 16481 1988
rect 18505 -1988 18539 1988
rect 20563 -1988 20597 1988
rect 22621 -1988 22655 1988
rect 24679 -1988 24713 1988
rect 26737 -1988 26771 1988
rect 28795 -1988 28829 1988
rect 30853 -1988 30887 1988
rect 32911 -1988 32945 1988
<< psubdiff >>
rect -33059 2140 -32963 2174
rect 32963 2140 33059 2174
rect -33059 2078 -33025 2140
rect 33025 2078 33059 2140
rect -33059 -2140 -33025 -2078
rect 33025 -2140 33059 -2078
rect -33059 -2174 -32963 -2140
rect 32963 -2174 33059 -2140
<< psubdiffcont >>
rect -32963 2140 32963 2174
rect -33059 -2078 -33025 2078
rect 33025 -2078 33059 2078
rect -32963 -2174 32963 -2140
<< poly >>
rect -32899 2072 -30899 2088
rect -32899 2038 -32883 2072
rect -30915 2038 -30899 2072
rect -32899 2000 -30899 2038
rect -30841 2072 -28841 2088
rect -30841 2038 -30825 2072
rect -28857 2038 -28841 2072
rect -30841 2000 -28841 2038
rect -28783 2072 -26783 2088
rect -28783 2038 -28767 2072
rect -26799 2038 -26783 2072
rect -28783 2000 -26783 2038
rect -26725 2072 -24725 2088
rect -26725 2038 -26709 2072
rect -24741 2038 -24725 2072
rect -26725 2000 -24725 2038
rect -24667 2072 -22667 2088
rect -24667 2038 -24651 2072
rect -22683 2038 -22667 2072
rect -24667 2000 -22667 2038
rect -22609 2072 -20609 2088
rect -22609 2038 -22593 2072
rect -20625 2038 -20609 2072
rect -22609 2000 -20609 2038
rect -20551 2072 -18551 2088
rect -20551 2038 -20535 2072
rect -18567 2038 -18551 2072
rect -20551 2000 -18551 2038
rect -18493 2072 -16493 2088
rect -18493 2038 -18477 2072
rect -16509 2038 -16493 2072
rect -18493 2000 -16493 2038
rect -16435 2072 -14435 2088
rect -16435 2038 -16419 2072
rect -14451 2038 -14435 2072
rect -16435 2000 -14435 2038
rect -14377 2072 -12377 2088
rect -14377 2038 -14361 2072
rect -12393 2038 -12377 2072
rect -14377 2000 -12377 2038
rect -12319 2072 -10319 2088
rect -12319 2038 -12303 2072
rect -10335 2038 -10319 2072
rect -12319 2000 -10319 2038
rect -10261 2072 -8261 2088
rect -10261 2038 -10245 2072
rect -8277 2038 -8261 2072
rect -10261 2000 -8261 2038
rect -8203 2072 -6203 2088
rect -8203 2038 -8187 2072
rect -6219 2038 -6203 2072
rect -8203 2000 -6203 2038
rect -6145 2072 -4145 2088
rect -6145 2038 -6129 2072
rect -4161 2038 -4145 2072
rect -6145 2000 -4145 2038
rect -4087 2072 -2087 2088
rect -4087 2038 -4071 2072
rect -2103 2038 -2087 2072
rect -4087 2000 -2087 2038
rect -2029 2072 -29 2088
rect -2029 2038 -2013 2072
rect -45 2038 -29 2072
rect -2029 2000 -29 2038
rect 29 2072 2029 2088
rect 29 2038 45 2072
rect 2013 2038 2029 2072
rect 29 2000 2029 2038
rect 2087 2072 4087 2088
rect 2087 2038 2103 2072
rect 4071 2038 4087 2072
rect 2087 2000 4087 2038
rect 4145 2072 6145 2088
rect 4145 2038 4161 2072
rect 6129 2038 6145 2072
rect 4145 2000 6145 2038
rect 6203 2072 8203 2088
rect 6203 2038 6219 2072
rect 8187 2038 8203 2072
rect 6203 2000 8203 2038
rect 8261 2072 10261 2088
rect 8261 2038 8277 2072
rect 10245 2038 10261 2072
rect 8261 2000 10261 2038
rect 10319 2072 12319 2088
rect 10319 2038 10335 2072
rect 12303 2038 12319 2072
rect 10319 2000 12319 2038
rect 12377 2072 14377 2088
rect 12377 2038 12393 2072
rect 14361 2038 14377 2072
rect 12377 2000 14377 2038
rect 14435 2072 16435 2088
rect 14435 2038 14451 2072
rect 16419 2038 16435 2072
rect 14435 2000 16435 2038
rect 16493 2072 18493 2088
rect 16493 2038 16509 2072
rect 18477 2038 18493 2072
rect 16493 2000 18493 2038
rect 18551 2072 20551 2088
rect 18551 2038 18567 2072
rect 20535 2038 20551 2072
rect 18551 2000 20551 2038
rect 20609 2072 22609 2088
rect 20609 2038 20625 2072
rect 22593 2038 22609 2072
rect 20609 2000 22609 2038
rect 22667 2072 24667 2088
rect 22667 2038 22683 2072
rect 24651 2038 24667 2072
rect 22667 2000 24667 2038
rect 24725 2072 26725 2088
rect 24725 2038 24741 2072
rect 26709 2038 26725 2072
rect 24725 2000 26725 2038
rect 26783 2072 28783 2088
rect 26783 2038 26799 2072
rect 28767 2038 28783 2072
rect 26783 2000 28783 2038
rect 28841 2072 30841 2088
rect 28841 2038 28857 2072
rect 30825 2038 30841 2072
rect 28841 2000 30841 2038
rect 30899 2072 32899 2088
rect 30899 2038 30915 2072
rect 32883 2038 32899 2072
rect 30899 2000 32899 2038
rect -32899 -2038 -30899 -2000
rect -32899 -2072 -32883 -2038
rect -30915 -2072 -30899 -2038
rect -32899 -2088 -30899 -2072
rect -30841 -2038 -28841 -2000
rect -30841 -2072 -30825 -2038
rect -28857 -2072 -28841 -2038
rect -30841 -2088 -28841 -2072
rect -28783 -2038 -26783 -2000
rect -28783 -2072 -28767 -2038
rect -26799 -2072 -26783 -2038
rect -28783 -2088 -26783 -2072
rect -26725 -2038 -24725 -2000
rect -26725 -2072 -26709 -2038
rect -24741 -2072 -24725 -2038
rect -26725 -2088 -24725 -2072
rect -24667 -2038 -22667 -2000
rect -24667 -2072 -24651 -2038
rect -22683 -2072 -22667 -2038
rect -24667 -2088 -22667 -2072
rect -22609 -2038 -20609 -2000
rect -22609 -2072 -22593 -2038
rect -20625 -2072 -20609 -2038
rect -22609 -2088 -20609 -2072
rect -20551 -2038 -18551 -2000
rect -20551 -2072 -20535 -2038
rect -18567 -2072 -18551 -2038
rect -20551 -2088 -18551 -2072
rect -18493 -2038 -16493 -2000
rect -18493 -2072 -18477 -2038
rect -16509 -2072 -16493 -2038
rect -18493 -2088 -16493 -2072
rect -16435 -2038 -14435 -2000
rect -16435 -2072 -16419 -2038
rect -14451 -2072 -14435 -2038
rect -16435 -2088 -14435 -2072
rect -14377 -2038 -12377 -2000
rect -14377 -2072 -14361 -2038
rect -12393 -2072 -12377 -2038
rect -14377 -2088 -12377 -2072
rect -12319 -2038 -10319 -2000
rect -12319 -2072 -12303 -2038
rect -10335 -2072 -10319 -2038
rect -12319 -2088 -10319 -2072
rect -10261 -2038 -8261 -2000
rect -10261 -2072 -10245 -2038
rect -8277 -2072 -8261 -2038
rect -10261 -2088 -8261 -2072
rect -8203 -2038 -6203 -2000
rect -8203 -2072 -8187 -2038
rect -6219 -2072 -6203 -2038
rect -8203 -2088 -6203 -2072
rect -6145 -2038 -4145 -2000
rect -6145 -2072 -6129 -2038
rect -4161 -2072 -4145 -2038
rect -6145 -2088 -4145 -2072
rect -4087 -2038 -2087 -2000
rect -4087 -2072 -4071 -2038
rect -2103 -2072 -2087 -2038
rect -4087 -2088 -2087 -2072
rect -2029 -2038 -29 -2000
rect -2029 -2072 -2013 -2038
rect -45 -2072 -29 -2038
rect -2029 -2088 -29 -2072
rect 29 -2038 2029 -2000
rect 29 -2072 45 -2038
rect 2013 -2072 2029 -2038
rect 29 -2088 2029 -2072
rect 2087 -2038 4087 -2000
rect 2087 -2072 2103 -2038
rect 4071 -2072 4087 -2038
rect 2087 -2088 4087 -2072
rect 4145 -2038 6145 -2000
rect 4145 -2072 4161 -2038
rect 6129 -2072 6145 -2038
rect 4145 -2088 6145 -2072
rect 6203 -2038 8203 -2000
rect 6203 -2072 6219 -2038
rect 8187 -2072 8203 -2038
rect 6203 -2088 8203 -2072
rect 8261 -2038 10261 -2000
rect 8261 -2072 8277 -2038
rect 10245 -2072 10261 -2038
rect 8261 -2088 10261 -2072
rect 10319 -2038 12319 -2000
rect 10319 -2072 10335 -2038
rect 12303 -2072 12319 -2038
rect 10319 -2088 12319 -2072
rect 12377 -2038 14377 -2000
rect 12377 -2072 12393 -2038
rect 14361 -2072 14377 -2038
rect 12377 -2088 14377 -2072
rect 14435 -2038 16435 -2000
rect 14435 -2072 14451 -2038
rect 16419 -2072 16435 -2038
rect 14435 -2088 16435 -2072
rect 16493 -2038 18493 -2000
rect 16493 -2072 16509 -2038
rect 18477 -2072 18493 -2038
rect 16493 -2088 18493 -2072
rect 18551 -2038 20551 -2000
rect 18551 -2072 18567 -2038
rect 20535 -2072 20551 -2038
rect 18551 -2088 20551 -2072
rect 20609 -2038 22609 -2000
rect 20609 -2072 20625 -2038
rect 22593 -2072 22609 -2038
rect 20609 -2088 22609 -2072
rect 22667 -2038 24667 -2000
rect 22667 -2072 22683 -2038
rect 24651 -2072 24667 -2038
rect 22667 -2088 24667 -2072
rect 24725 -2038 26725 -2000
rect 24725 -2072 24741 -2038
rect 26709 -2072 26725 -2038
rect 24725 -2088 26725 -2072
rect 26783 -2038 28783 -2000
rect 26783 -2072 26799 -2038
rect 28767 -2072 28783 -2038
rect 26783 -2088 28783 -2072
rect 28841 -2038 30841 -2000
rect 28841 -2072 28857 -2038
rect 30825 -2072 30841 -2038
rect 28841 -2088 30841 -2072
rect 30899 -2038 32899 -2000
rect 30899 -2072 30915 -2038
rect 32883 -2072 32899 -2038
rect 30899 -2088 32899 -2072
<< polycont >>
rect -32883 2038 -30915 2072
rect -30825 2038 -28857 2072
rect -28767 2038 -26799 2072
rect -26709 2038 -24741 2072
rect -24651 2038 -22683 2072
rect -22593 2038 -20625 2072
rect -20535 2038 -18567 2072
rect -18477 2038 -16509 2072
rect -16419 2038 -14451 2072
rect -14361 2038 -12393 2072
rect -12303 2038 -10335 2072
rect -10245 2038 -8277 2072
rect -8187 2038 -6219 2072
rect -6129 2038 -4161 2072
rect -4071 2038 -2103 2072
rect -2013 2038 -45 2072
rect 45 2038 2013 2072
rect 2103 2038 4071 2072
rect 4161 2038 6129 2072
rect 6219 2038 8187 2072
rect 8277 2038 10245 2072
rect 10335 2038 12303 2072
rect 12393 2038 14361 2072
rect 14451 2038 16419 2072
rect 16509 2038 18477 2072
rect 18567 2038 20535 2072
rect 20625 2038 22593 2072
rect 22683 2038 24651 2072
rect 24741 2038 26709 2072
rect 26799 2038 28767 2072
rect 28857 2038 30825 2072
rect 30915 2038 32883 2072
rect -32883 -2072 -30915 -2038
rect -30825 -2072 -28857 -2038
rect -28767 -2072 -26799 -2038
rect -26709 -2072 -24741 -2038
rect -24651 -2072 -22683 -2038
rect -22593 -2072 -20625 -2038
rect -20535 -2072 -18567 -2038
rect -18477 -2072 -16509 -2038
rect -16419 -2072 -14451 -2038
rect -14361 -2072 -12393 -2038
rect -12303 -2072 -10335 -2038
rect -10245 -2072 -8277 -2038
rect -8187 -2072 -6219 -2038
rect -6129 -2072 -4161 -2038
rect -4071 -2072 -2103 -2038
rect -2013 -2072 -45 -2038
rect 45 -2072 2013 -2038
rect 2103 -2072 4071 -2038
rect 4161 -2072 6129 -2038
rect 6219 -2072 8187 -2038
rect 8277 -2072 10245 -2038
rect 10335 -2072 12303 -2038
rect 12393 -2072 14361 -2038
rect 14451 -2072 16419 -2038
rect 16509 -2072 18477 -2038
rect 18567 -2072 20535 -2038
rect 20625 -2072 22593 -2038
rect 22683 -2072 24651 -2038
rect 24741 -2072 26709 -2038
rect 26799 -2072 28767 -2038
rect 28857 -2072 30825 -2038
rect 30915 -2072 32883 -2038
<< locali >>
rect -33059 2140 -32963 2174
rect 32963 2140 33059 2174
rect -33059 2078 -33025 2140
rect 33025 2078 33059 2140
rect -32899 2038 -32883 2072
rect -30915 2038 -30899 2072
rect -30841 2038 -30825 2072
rect -28857 2038 -28841 2072
rect -28783 2038 -28767 2072
rect -26799 2038 -26783 2072
rect -26725 2038 -26709 2072
rect -24741 2038 -24725 2072
rect -24667 2038 -24651 2072
rect -22683 2038 -22667 2072
rect -22609 2038 -22593 2072
rect -20625 2038 -20609 2072
rect -20551 2038 -20535 2072
rect -18567 2038 -18551 2072
rect -18493 2038 -18477 2072
rect -16509 2038 -16493 2072
rect -16435 2038 -16419 2072
rect -14451 2038 -14435 2072
rect -14377 2038 -14361 2072
rect -12393 2038 -12377 2072
rect -12319 2038 -12303 2072
rect -10335 2038 -10319 2072
rect -10261 2038 -10245 2072
rect -8277 2038 -8261 2072
rect -8203 2038 -8187 2072
rect -6219 2038 -6203 2072
rect -6145 2038 -6129 2072
rect -4161 2038 -4145 2072
rect -4087 2038 -4071 2072
rect -2103 2038 -2087 2072
rect -2029 2038 -2013 2072
rect -45 2038 -29 2072
rect 29 2038 45 2072
rect 2013 2038 2029 2072
rect 2087 2038 2103 2072
rect 4071 2038 4087 2072
rect 4145 2038 4161 2072
rect 6129 2038 6145 2072
rect 6203 2038 6219 2072
rect 8187 2038 8203 2072
rect 8261 2038 8277 2072
rect 10245 2038 10261 2072
rect 10319 2038 10335 2072
rect 12303 2038 12319 2072
rect 12377 2038 12393 2072
rect 14361 2038 14377 2072
rect 14435 2038 14451 2072
rect 16419 2038 16435 2072
rect 16493 2038 16509 2072
rect 18477 2038 18493 2072
rect 18551 2038 18567 2072
rect 20535 2038 20551 2072
rect 20609 2038 20625 2072
rect 22593 2038 22609 2072
rect 22667 2038 22683 2072
rect 24651 2038 24667 2072
rect 24725 2038 24741 2072
rect 26709 2038 26725 2072
rect 26783 2038 26799 2072
rect 28767 2038 28783 2072
rect 28841 2038 28857 2072
rect 30825 2038 30841 2072
rect 30899 2038 30915 2072
rect 32883 2038 32899 2072
rect -32945 1988 -32911 2004
rect -32945 -2004 -32911 -1988
rect -30887 1988 -30853 2004
rect -30887 -2004 -30853 -1988
rect -28829 1988 -28795 2004
rect -28829 -2004 -28795 -1988
rect -26771 1988 -26737 2004
rect -26771 -2004 -26737 -1988
rect -24713 1988 -24679 2004
rect -24713 -2004 -24679 -1988
rect -22655 1988 -22621 2004
rect -22655 -2004 -22621 -1988
rect -20597 1988 -20563 2004
rect -20597 -2004 -20563 -1988
rect -18539 1988 -18505 2004
rect -18539 -2004 -18505 -1988
rect -16481 1988 -16447 2004
rect -16481 -2004 -16447 -1988
rect -14423 1988 -14389 2004
rect -14423 -2004 -14389 -1988
rect -12365 1988 -12331 2004
rect -12365 -2004 -12331 -1988
rect -10307 1988 -10273 2004
rect -10307 -2004 -10273 -1988
rect -8249 1988 -8215 2004
rect -8249 -2004 -8215 -1988
rect -6191 1988 -6157 2004
rect -6191 -2004 -6157 -1988
rect -4133 1988 -4099 2004
rect -4133 -2004 -4099 -1988
rect -2075 1988 -2041 2004
rect -2075 -2004 -2041 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 2041 1988 2075 2004
rect 2041 -2004 2075 -1988
rect 4099 1988 4133 2004
rect 4099 -2004 4133 -1988
rect 6157 1988 6191 2004
rect 6157 -2004 6191 -1988
rect 8215 1988 8249 2004
rect 8215 -2004 8249 -1988
rect 10273 1988 10307 2004
rect 10273 -2004 10307 -1988
rect 12331 1988 12365 2004
rect 12331 -2004 12365 -1988
rect 14389 1988 14423 2004
rect 14389 -2004 14423 -1988
rect 16447 1988 16481 2004
rect 16447 -2004 16481 -1988
rect 18505 1988 18539 2004
rect 18505 -2004 18539 -1988
rect 20563 1988 20597 2004
rect 20563 -2004 20597 -1988
rect 22621 1988 22655 2004
rect 22621 -2004 22655 -1988
rect 24679 1988 24713 2004
rect 24679 -2004 24713 -1988
rect 26737 1988 26771 2004
rect 26737 -2004 26771 -1988
rect 28795 1988 28829 2004
rect 28795 -2004 28829 -1988
rect 30853 1988 30887 2004
rect 30853 -2004 30887 -1988
rect 32911 1988 32945 2004
rect 32911 -2004 32945 -1988
rect -32899 -2072 -32883 -2038
rect -30915 -2072 -30899 -2038
rect -30841 -2072 -30825 -2038
rect -28857 -2072 -28841 -2038
rect -28783 -2072 -28767 -2038
rect -26799 -2072 -26783 -2038
rect -26725 -2072 -26709 -2038
rect -24741 -2072 -24725 -2038
rect -24667 -2072 -24651 -2038
rect -22683 -2072 -22667 -2038
rect -22609 -2072 -22593 -2038
rect -20625 -2072 -20609 -2038
rect -20551 -2072 -20535 -2038
rect -18567 -2072 -18551 -2038
rect -18493 -2072 -18477 -2038
rect -16509 -2072 -16493 -2038
rect -16435 -2072 -16419 -2038
rect -14451 -2072 -14435 -2038
rect -14377 -2072 -14361 -2038
rect -12393 -2072 -12377 -2038
rect -12319 -2072 -12303 -2038
rect -10335 -2072 -10319 -2038
rect -10261 -2072 -10245 -2038
rect -8277 -2072 -8261 -2038
rect -8203 -2072 -8187 -2038
rect -6219 -2072 -6203 -2038
rect -6145 -2072 -6129 -2038
rect -4161 -2072 -4145 -2038
rect -4087 -2072 -4071 -2038
rect -2103 -2072 -2087 -2038
rect -2029 -2072 -2013 -2038
rect -45 -2072 -29 -2038
rect 29 -2072 45 -2038
rect 2013 -2072 2029 -2038
rect 2087 -2072 2103 -2038
rect 4071 -2072 4087 -2038
rect 4145 -2072 4161 -2038
rect 6129 -2072 6145 -2038
rect 6203 -2072 6219 -2038
rect 8187 -2072 8203 -2038
rect 8261 -2072 8277 -2038
rect 10245 -2072 10261 -2038
rect 10319 -2072 10335 -2038
rect 12303 -2072 12319 -2038
rect 12377 -2072 12393 -2038
rect 14361 -2072 14377 -2038
rect 14435 -2072 14451 -2038
rect 16419 -2072 16435 -2038
rect 16493 -2072 16509 -2038
rect 18477 -2072 18493 -2038
rect 18551 -2072 18567 -2038
rect 20535 -2072 20551 -2038
rect 20609 -2072 20625 -2038
rect 22593 -2072 22609 -2038
rect 22667 -2072 22683 -2038
rect 24651 -2072 24667 -2038
rect 24725 -2072 24741 -2038
rect 26709 -2072 26725 -2038
rect 26783 -2072 26799 -2038
rect 28767 -2072 28783 -2038
rect 28841 -2072 28857 -2038
rect 30825 -2072 30841 -2038
rect 30899 -2072 30915 -2038
rect 32883 -2072 32899 -2038
rect -33059 -2140 -33025 -2078
rect 33025 -2140 33059 -2078
rect -33059 -2174 -32963 -2140
rect 32963 -2174 33059 -2140
<< viali >>
rect -32883 2038 -30915 2072
rect -30825 2038 -28857 2072
rect -28767 2038 -26799 2072
rect -26709 2038 -24741 2072
rect -24651 2038 -22683 2072
rect -22593 2038 -20625 2072
rect -20535 2038 -18567 2072
rect -18477 2038 -16509 2072
rect -16419 2038 -14451 2072
rect -14361 2038 -12393 2072
rect -12303 2038 -10335 2072
rect -10245 2038 -8277 2072
rect -8187 2038 -6219 2072
rect -6129 2038 -4161 2072
rect -4071 2038 -2103 2072
rect -2013 2038 -45 2072
rect 45 2038 2013 2072
rect 2103 2038 4071 2072
rect 4161 2038 6129 2072
rect 6219 2038 8187 2072
rect 8277 2038 10245 2072
rect 10335 2038 12303 2072
rect 12393 2038 14361 2072
rect 14451 2038 16419 2072
rect 16509 2038 18477 2072
rect 18567 2038 20535 2072
rect 20625 2038 22593 2072
rect 22683 2038 24651 2072
rect 24741 2038 26709 2072
rect 26799 2038 28767 2072
rect 28857 2038 30825 2072
rect 30915 2038 32883 2072
rect -32945 -1988 -32911 1988
rect -30887 -1988 -30853 1988
rect -28829 -1988 -28795 1988
rect -26771 -1988 -26737 1988
rect -24713 -1988 -24679 1988
rect -22655 -1988 -22621 1988
rect -20597 -1988 -20563 1988
rect -18539 -1988 -18505 1988
rect -16481 -1988 -16447 1988
rect -14423 -1988 -14389 1988
rect -12365 -1988 -12331 1988
rect -10307 -1988 -10273 1988
rect -8249 -1988 -8215 1988
rect -6191 -1988 -6157 1988
rect -4133 -1988 -4099 1988
rect -2075 -1988 -2041 1988
rect -17 -1988 17 1988
rect 2041 -1988 2075 1988
rect 4099 -1988 4133 1988
rect 6157 -1988 6191 1988
rect 8215 -1988 8249 1988
rect 10273 -1988 10307 1988
rect 12331 -1988 12365 1988
rect 14389 -1988 14423 1988
rect 16447 -1988 16481 1988
rect 18505 -1988 18539 1988
rect 20563 -1988 20597 1988
rect 22621 -1988 22655 1988
rect 24679 -1988 24713 1988
rect 26737 -1988 26771 1988
rect 28795 -1988 28829 1988
rect 30853 -1988 30887 1988
rect 32911 -1988 32945 1988
rect -32883 -2072 -30915 -2038
rect -30825 -2072 -28857 -2038
rect -28767 -2072 -26799 -2038
rect -26709 -2072 -24741 -2038
rect -24651 -2072 -22683 -2038
rect -22593 -2072 -20625 -2038
rect -20535 -2072 -18567 -2038
rect -18477 -2072 -16509 -2038
rect -16419 -2072 -14451 -2038
rect -14361 -2072 -12393 -2038
rect -12303 -2072 -10335 -2038
rect -10245 -2072 -8277 -2038
rect -8187 -2072 -6219 -2038
rect -6129 -2072 -4161 -2038
rect -4071 -2072 -2103 -2038
rect -2013 -2072 -45 -2038
rect 45 -2072 2013 -2038
rect 2103 -2072 4071 -2038
rect 4161 -2072 6129 -2038
rect 6219 -2072 8187 -2038
rect 8277 -2072 10245 -2038
rect 10335 -2072 12303 -2038
rect 12393 -2072 14361 -2038
rect 14451 -2072 16419 -2038
rect 16509 -2072 18477 -2038
rect 18567 -2072 20535 -2038
rect 20625 -2072 22593 -2038
rect 22683 -2072 24651 -2038
rect 24741 -2072 26709 -2038
rect 26799 -2072 28767 -2038
rect 28857 -2072 30825 -2038
rect 30915 -2072 32883 -2038
<< metal1 >>
rect -32895 2072 -30903 2078
rect -32895 2038 -32883 2072
rect -30915 2038 -30903 2072
rect -32895 2032 -30903 2038
rect -30837 2072 -28845 2078
rect -30837 2038 -30825 2072
rect -28857 2038 -28845 2072
rect -30837 2032 -28845 2038
rect -28779 2072 -26787 2078
rect -28779 2038 -28767 2072
rect -26799 2038 -26787 2072
rect -28779 2032 -26787 2038
rect -26721 2072 -24729 2078
rect -26721 2038 -26709 2072
rect -24741 2038 -24729 2072
rect -26721 2032 -24729 2038
rect -24663 2072 -22671 2078
rect -24663 2038 -24651 2072
rect -22683 2038 -22671 2072
rect -24663 2032 -22671 2038
rect -22605 2072 -20613 2078
rect -22605 2038 -22593 2072
rect -20625 2038 -20613 2072
rect -22605 2032 -20613 2038
rect -20547 2072 -18555 2078
rect -20547 2038 -20535 2072
rect -18567 2038 -18555 2072
rect -20547 2032 -18555 2038
rect -18489 2072 -16497 2078
rect -18489 2038 -18477 2072
rect -16509 2038 -16497 2072
rect -18489 2032 -16497 2038
rect -16431 2072 -14439 2078
rect -16431 2038 -16419 2072
rect -14451 2038 -14439 2072
rect -16431 2032 -14439 2038
rect -14373 2072 -12381 2078
rect -14373 2038 -14361 2072
rect -12393 2038 -12381 2072
rect -14373 2032 -12381 2038
rect -12315 2072 -10323 2078
rect -12315 2038 -12303 2072
rect -10335 2038 -10323 2072
rect -12315 2032 -10323 2038
rect -10257 2072 -8265 2078
rect -10257 2038 -10245 2072
rect -8277 2038 -8265 2072
rect -10257 2032 -8265 2038
rect -8199 2072 -6207 2078
rect -8199 2038 -8187 2072
rect -6219 2038 -6207 2072
rect -8199 2032 -6207 2038
rect -6141 2072 -4149 2078
rect -6141 2038 -6129 2072
rect -4161 2038 -4149 2072
rect -6141 2032 -4149 2038
rect -4083 2072 -2091 2078
rect -4083 2038 -4071 2072
rect -2103 2038 -2091 2072
rect -4083 2032 -2091 2038
rect -2025 2072 -33 2078
rect -2025 2038 -2013 2072
rect -45 2038 -33 2072
rect -2025 2032 -33 2038
rect 33 2072 2025 2078
rect 33 2038 45 2072
rect 2013 2038 2025 2072
rect 33 2032 2025 2038
rect 2091 2072 4083 2078
rect 2091 2038 2103 2072
rect 4071 2038 4083 2072
rect 2091 2032 4083 2038
rect 4149 2072 6141 2078
rect 4149 2038 4161 2072
rect 6129 2038 6141 2072
rect 4149 2032 6141 2038
rect 6207 2072 8199 2078
rect 6207 2038 6219 2072
rect 8187 2038 8199 2072
rect 6207 2032 8199 2038
rect 8265 2072 10257 2078
rect 8265 2038 8277 2072
rect 10245 2038 10257 2072
rect 8265 2032 10257 2038
rect 10323 2072 12315 2078
rect 10323 2038 10335 2072
rect 12303 2038 12315 2072
rect 10323 2032 12315 2038
rect 12381 2072 14373 2078
rect 12381 2038 12393 2072
rect 14361 2038 14373 2072
rect 12381 2032 14373 2038
rect 14439 2072 16431 2078
rect 14439 2038 14451 2072
rect 16419 2038 16431 2072
rect 14439 2032 16431 2038
rect 16497 2072 18489 2078
rect 16497 2038 16509 2072
rect 18477 2038 18489 2072
rect 16497 2032 18489 2038
rect 18555 2072 20547 2078
rect 18555 2038 18567 2072
rect 20535 2038 20547 2072
rect 18555 2032 20547 2038
rect 20613 2072 22605 2078
rect 20613 2038 20625 2072
rect 22593 2038 22605 2072
rect 20613 2032 22605 2038
rect 22671 2072 24663 2078
rect 22671 2038 22683 2072
rect 24651 2038 24663 2072
rect 22671 2032 24663 2038
rect 24729 2072 26721 2078
rect 24729 2038 24741 2072
rect 26709 2038 26721 2072
rect 24729 2032 26721 2038
rect 26787 2072 28779 2078
rect 26787 2038 26799 2072
rect 28767 2038 28779 2072
rect 26787 2032 28779 2038
rect 28845 2072 30837 2078
rect 28845 2038 28857 2072
rect 30825 2038 30837 2072
rect 28845 2032 30837 2038
rect 30903 2072 32895 2078
rect 30903 2038 30915 2072
rect 32883 2038 32895 2072
rect 30903 2032 32895 2038
rect -32951 1988 -32905 2000
rect -32951 -1988 -32945 1988
rect -32911 -1988 -32905 1988
rect -32951 -2000 -32905 -1988
rect -30893 1988 -30847 2000
rect -30893 -1988 -30887 1988
rect -30853 -1988 -30847 1988
rect -30893 -2000 -30847 -1988
rect -28835 1988 -28789 2000
rect -28835 -1988 -28829 1988
rect -28795 -1988 -28789 1988
rect -28835 -2000 -28789 -1988
rect -26777 1988 -26731 2000
rect -26777 -1988 -26771 1988
rect -26737 -1988 -26731 1988
rect -26777 -2000 -26731 -1988
rect -24719 1988 -24673 2000
rect -24719 -1988 -24713 1988
rect -24679 -1988 -24673 1988
rect -24719 -2000 -24673 -1988
rect -22661 1988 -22615 2000
rect -22661 -1988 -22655 1988
rect -22621 -1988 -22615 1988
rect -22661 -2000 -22615 -1988
rect -20603 1988 -20557 2000
rect -20603 -1988 -20597 1988
rect -20563 -1988 -20557 1988
rect -20603 -2000 -20557 -1988
rect -18545 1988 -18499 2000
rect -18545 -1988 -18539 1988
rect -18505 -1988 -18499 1988
rect -18545 -2000 -18499 -1988
rect -16487 1988 -16441 2000
rect -16487 -1988 -16481 1988
rect -16447 -1988 -16441 1988
rect -16487 -2000 -16441 -1988
rect -14429 1988 -14383 2000
rect -14429 -1988 -14423 1988
rect -14389 -1988 -14383 1988
rect -14429 -2000 -14383 -1988
rect -12371 1988 -12325 2000
rect -12371 -1988 -12365 1988
rect -12331 -1988 -12325 1988
rect -12371 -2000 -12325 -1988
rect -10313 1988 -10267 2000
rect -10313 -1988 -10307 1988
rect -10273 -1988 -10267 1988
rect -10313 -2000 -10267 -1988
rect -8255 1988 -8209 2000
rect -8255 -1988 -8249 1988
rect -8215 -1988 -8209 1988
rect -8255 -2000 -8209 -1988
rect -6197 1988 -6151 2000
rect -6197 -1988 -6191 1988
rect -6157 -1988 -6151 1988
rect -6197 -2000 -6151 -1988
rect -4139 1988 -4093 2000
rect -4139 -1988 -4133 1988
rect -4099 -1988 -4093 1988
rect -4139 -2000 -4093 -1988
rect -2081 1988 -2035 2000
rect -2081 -1988 -2075 1988
rect -2041 -1988 -2035 1988
rect -2081 -2000 -2035 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 2035 1988 2081 2000
rect 2035 -1988 2041 1988
rect 2075 -1988 2081 1988
rect 2035 -2000 2081 -1988
rect 4093 1988 4139 2000
rect 4093 -1988 4099 1988
rect 4133 -1988 4139 1988
rect 4093 -2000 4139 -1988
rect 6151 1988 6197 2000
rect 6151 -1988 6157 1988
rect 6191 -1988 6197 1988
rect 6151 -2000 6197 -1988
rect 8209 1988 8255 2000
rect 8209 -1988 8215 1988
rect 8249 -1988 8255 1988
rect 8209 -2000 8255 -1988
rect 10267 1988 10313 2000
rect 10267 -1988 10273 1988
rect 10307 -1988 10313 1988
rect 10267 -2000 10313 -1988
rect 12325 1988 12371 2000
rect 12325 -1988 12331 1988
rect 12365 -1988 12371 1988
rect 12325 -2000 12371 -1988
rect 14383 1988 14429 2000
rect 14383 -1988 14389 1988
rect 14423 -1988 14429 1988
rect 14383 -2000 14429 -1988
rect 16441 1988 16487 2000
rect 16441 -1988 16447 1988
rect 16481 -1988 16487 1988
rect 16441 -2000 16487 -1988
rect 18499 1988 18545 2000
rect 18499 -1988 18505 1988
rect 18539 -1988 18545 1988
rect 18499 -2000 18545 -1988
rect 20557 1988 20603 2000
rect 20557 -1988 20563 1988
rect 20597 -1988 20603 1988
rect 20557 -2000 20603 -1988
rect 22615 1988 22661 2000
rect 22615 -1988 22621 1988
rect 22655 -1988 22661 1988
rect 22615 -2000 22661 -1988
rect 24673 1988 24719 2000
rect 24673 -1988 24679 1988
rect 24713 -1988 24719 1988
rect 24673 -2000 24719 -1988
rect 26731 1988 26777 2000
rect 26731 -1988 26737 1988
rect 26771 -1988 26777 1988
rect 26731 -2000 26777 -1988
rect 28789 1988 28835 2000
rect 28789 -1988 28795 1988
rect 28829 -1988 28835 1988
rect 28789 -2000 28835 -1988
rect 30847 1988 30893 2000
rect 30847 -1988 30853 1988
rect 30887 -1988 30893 1988
rect 30847 -2000 30893 -1988
rect 32905 1988 32951 2000
rect 32905 -1988 32911 1988
rect 32945 -1988 32951 1988
rect 32905 -2000 32951 -1988
rect -32895 -2038 -30903 -2032
rect -32895 -2072 -32883 -2038
rect -30915 -2072 -30903 -2038
rect -32895 -2078 -30903 -2072
rect -30837 -2038 -28845 -2032
rect -30837 -2072 -30825 -2038
rect -28857 -2072 -28845 -2038
rect -30837 -2078 -28845 -2072
rect -28779 -2038 -26787 -2032
rect -28779 -2072 -28767 -2038
rect -26799 -2072 -26787 -2038
rect -28779 -2078 -26787 -2072
rect -26721 -2038 -24729 -2032
rect -26721 -2072 -26709 -2038
rect -24741 -2072 -24729 -2038
rect -26721 -2078 -24729 -2072
rect -24663 -2038 -22671 -2032
rect -24663 -2072 -24651 -2038
rect -22683 -2072 -22671 -2038
rect -24663 -2078 -22671 -2072
rect -22605 -2038 -20613 -2032
rect -22605 -2072 -22593 -2038
rect -20625 -2072 -20613 -2038
rect -22605 -2078 -20613 -2072
rect -20547 -2038 -18555 -2032
rect -20547 -2072 -20535 -2038
rect -18567 -2072 -18555 -2038
rect -20547 -2078 -18555 -2072
rect -18489 -2038 -16497 -2032
rect -18489 -2072 -18477 -2038
rect -16509 -2072 -16497 -2038
rect -18489 -2078 -16497 -2072
rect -16431 -2038 -14439 -2032
rect -16431 -2072 -16419 -2038
rect -14451 -2072 -14439 -2038
rect -16431 -2078 -14439 -2072
rect -14373 -2038 -12381 -2032
rect -14373 -2072 -14361 -2038
rect -12393 -2072 -12381 -2038
rect -14373 -2078 -12381 -2072
rect -12315 -2038 -10323 -2032
rect -12315 -2072 -12303 -2038
rect -10335 -2072 -10323 -2038
rect -12315 -2078 -10323 -2072
rect -10257 -2038 -8265 -2032
rect -10257 -2072 -10245 -2038
rect -8277 -2072 -8265 -2038
rect -10257 -2078 -8265 -2072
rect -8199 -2038 -6207 -2032
rect -8199 -2072 -8187 -2038
rect -6219 -2072 -6207 -2038
rect -8199 -2078 -6207 -2072
rect -6141 -2038 -4149 -2032
rect -6141 -2072 -6129 -2038
rect -4161 -2072 -4149 -2038
rect -6141 -2078 -4149 -2072
rect -4083 -2038 -2091 -2032
rect -4083 -2072 -4071 -2038
rect -2103 -2072 -2091 -2038
rect -4083 -2078 -2091 -2072
rect -2025 -2038 -33 -2032
rect -2025 -2072 -2013 -2038
rect -45 -2072 -33 -2038
rect -2025 -2078 -33 -2072
rect 33 -2038 2025 -2032
rect 33 -2072 45 -2038
rect 2013 -2072 2025 -2038
rect 33 -2078 2025 -2072
rect 2091 -2038 4083 -2032
rect 2091 -2072 2103 -2038
rect 4071 -2072 4083 -2038
rect 2091 -2078 4083 -2072
rect 4149 -2038 6141 -2032
rect 4149 -2072 4161 -2038
rect 6129 -2072 6141 -2038
rect 4149 -2078 6141 -2072
rect 6207 -2038 8199 -2032
rect 6207 -2072 6219 -2038
rect 8187 -2072 8199 -2038
rect 6207 -2078 8199 -2072
rect 8265 -2038 10257 -2032
rect 8265 -2072 8277 -2038
rect 10245 -2072 10257 -2038
rect 8265 -2078 10257 -2072
rect 10323 -2038 12315 -2032
rect 10323 -2072 10335 -2038
rect 12303 -2072 12315 -2038
rect 10323 -2078 12315 -2072
rect 12381 -2038 14373 -2032
rect 12381 -2072 12393 -2038
rect 14361 -2072 14373 -2038
rect 12381 -2078 14373 -2072
rect 14439 -2038 16431 -2032
rect 14439 -2072 14451 -2038
rect 16419 -2072 16431 -2038
rect 14439 -2078 16431 -2072
rect 16497 -2038 18489 -2032
rect 16497 -2072 16509 -2038
rect 18477 -2072 18489 -2038
rect 16497 -2078 18489 -2072
rect 18555 -2038 20547 -2032
rect 18555 -2072 18567 -2038
rect 20535 -2072 20547 -2038
rect 18555 -2078 20547 -2072
rect 20613 -2038 22605 -2032
rect 20613 -2072 20625 -2038
rect 22593 -2072 22605 -2038
rect 20613 -2078 22605 -2072
rect 22671 -2038 24663 -2032
rect 22671 -2072 22683 -2038
rect 24651 -2072 24663 -2038
rect 22671 -2078 24663 -2072
rect 24729 -2038 26721 -2032
rect 24729 -2072 24741 -2038
rect 26709 -2072 26721 -2038
rect 24729 -2078 26721 -2072
rect 26787 -2038 28779 -2032
rect 26787 -2072 26799 -2038
rect 28767 -2072 28779 -2038
rect 26787 -2078 28779 -2072
rect 28845 -2038 30837 -2032
rect 28845 -2072 28857 -2038
rect 30825 -2072 30837 -2038
rect 28845 -2078 30837 -2072
rect 30903 -2038 32895 -2032
rect 30903 -2072 30915 -2038
rect 32883 -2072 32895 -2038
rect 30903 -2078 32895 -2072
<< properties >>
string FIXED_BBOX -33042 -2157 33042 2157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20 l 10 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
