magic
tech sky130A
magscale 1 2
timestamp 1697806833
<< nwell >>
rect -3254 -4219 3254 4219
<< pmos >>
rect -3058 -4000 -1058 4000
rect -1000 -4000 1000 4000
rect 1058 -4000 3058 4000
<< pdiff >>
rect -3116 3988 -3058 4000
rect -3116 -3988 -3104 3988
rect -3070 -3988 -3058 3988
rect -3116 -4000 -3058 -3988
rect -1058 3988 -1000 4000
rect -1058 -3988 -1046 3988
rect -1012 -3988 -1000 3988
rect -1058 -4000 -1000 -3988
rect 1000 3988 1058 4000
rect 1000 -3988 1012 3988
rect 1046 -3988 1058 3988
rect 1000 -4000 1058 -3988
rect 3058 3988 3116 4000
rect 3058 -3988 3070 3988
rect 3104 -3988 3116 3988
rect 3058 -4000 3116 -3988
<< pdiffc >>
rect -3104 -3988 -3070 3988
rect -1046 -3988 -1012 3988
rect 1012 -3988 1046 3988
rect 3070 -3988 3104 3988
<< nsubdiff >>
rect -3218 4149 -3122 4183
rect 3122 4149 3218 4183
rect -3218 4087 -3184 4149
rect 3184 4087 3218 4149
rect -3218 -4149 -3184 -4087
rect 3184 -4149 3218 -4087
rect -3218 -4183 -3122 -4149
rect 3122 -4183 3218 -4149
<< nsubdiffcont >>
rect -3122 4149 3122 4183
rect -3218 -4087 -3184 4087
rect 3184 -4087 3218 4087
rect -3122 -4183 3122 -4149
<< poly >>
rect -3058 4081 -1058 4097
rect -3058 4047 -3042 4081
rect -1074 4047 -1058 4081
rect -3058 4000 -1058 4047
rect -1000 4081 1000 4097
rect -1000 4047 -984 4081
rect 984 4047 1000 4081
rect -1000 4000 1000 4047
rect 1058 4081 3058 4097
rect 1058 4047 1074 4081
rect 3042 4047 3058 4081
rect 1058 4000 3058 4047
rect -3058 -4047 -1058 -4000
rect -3058 -4081 -3042 -4047
rect -1074 -4081 -1058 -4047
rect -3058 -4097 -1058 -4081
rect -1000 -4047 1000 -4000
rect -1000 -4081 -984 -4047
rect 984 -4081 1000 -4047
rect -1000 -4097 1000 -4081
rect 1058 -4047 3058 -4000
rect 1058 -4081 1074 -4047
rect 3042 -4081 3058 -4047
rect 1058 -4097 3058 -4081
<< polycont >>
rect -3042 4047 -1074 4081
rect -984 4047 984 4081
rect 1074 4047 3042 4081
rect -3042 -4081 -1074 -4047
rect -984 -4081 984 -4047
rect 1074 -4081 3042 -4047
<< locali >>
rect -3218 4149 -3122 4183
rect 3122 4149 3218 4183
rect -3218 4087 -3184 4149
rect 3184 4087 3218 4149
rect -3058 4047 -3042 4081
rect -1074 4047 -1058 4081
rect -1000 4047 -984 4081
rect 984 4047 1000 4081
rect 1058 4047 1074 4081
rect 3042 4047 3058 4081
rect -3104 3988 -3070 4004
rect -3104 -4004 -3070 -3988
rect -1046 3988 -1012 4004
rect -1046 -4004 -1012 -3988
rect 1012 3988 1046 4004
rect 1012 -4004 1046 -3988
rect 3070 3988 3104 4004
rect 3070 -4004 3104 -3988
rect -3058 -4081 -3042 -4047
rect -1074 -4081 -1058 -4047
rect -1000 -4081 -984 -4047
rect 984 -4081 1000 -4047
rect 1058 -4081 1074 -4047
rect 3042 -4081 3058 -4047
rect -3218 -4149 -3184 -4087
rect 3184 -4149 3218 -4087
rect -3218 -4183 -3122 -4149
rect 3122 -4183 3218 -4149
<< viali >>
rect -3042 4047 -1074 4081
rect -984 4047 984 4081
rect 1074 4047 3042 4081
rect -3104 -3988 -3070 3988
rect -1046 -3988 -1012 3988
rect 1012 -3988 1046 3988
rect 3070 -3988 3104 3988
rect -3042 -4081 -1074 -4047
rect -984 -4081 984 -4047
rect 1074 -4081 3042 -4047
<< metal1 >>
rect -3054 4081 -1062 4087
rect -3054 4047 -3042 4081
rect -1074 4047 -1062 4081
rect -3054 4041 -1062 4047
rect -996 4081 996 4087
rect -996 4047 -984 4081
rect 984 4047 996 4081
rect -996 4041 996 4047
rect 1062 4081 3054 4087
rect 1062 4047 1074 4081
rect 3042 4047 3054 4081
rect 1062 4041 3054 4047
rect -3110 3988 -3064 4000
rect -3110 -3988 -3104 3988
rect -3070 -3988 -3064 3988
rect -3110 -4000 -3064 -3988
rect -1052 3988 -1006 4000
rect -1052 -3988 -1046 3988
rect -1012 -3988 -1006 3988
rect -1052 -4000 -1006 -3988
rect 1006 3988 1052 4000
rect 1006 -3988 1012 3988
rect 1046 -3988 1052 3988
rect 1006 -4000 1052 -3988
rect 3064 3988 3110 4000
rect 3064 -3988 3070 3988
rect 3104 -3988 3110 3988
rect 3064 -4000 3110 -3988
rect -3054 -4047 -1062 -4041
rect -3054 -4081 -3042 -4047
rect -1074 -4081 -1062 -4047
rect -3054 -4087 -1062 -4081
rect -996 -4047 996 -4041
rect -996 -4081 -984 -4047
rect 984 -4081 996 -4047
rect -996 -4087 996 -4081
rect 1062 -4047 3054 -4041
rect 1062 -4081 1074 -4047
rect 3042 -4081 3054 -4047
rect 1062 -4087 3054 -4081
<< properties >>
string FIXED_BBOX -3201 -4166 3201 4166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 40 l 10 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
