magic
tech sky130A
magscale 1 2
timestamp 1697785254
<< locali >>
rect -8500 17500 -8000 18700
rect -9700 17000 -8000 17500
rect -8500 16950 -8000 17000
rect -7950 16950 -7450 18700
rect -9700 16450 -7450 16950
rect -7950 16400 -7450 16450
rect -7400 16400 -6900 18700
rect -9700 15900 -6900 16400
rect -7400 15850 -6900 15900
rect -6850 15850 -6350 18700
rect -9700 15350 -6350 15850
rect -6850 15300 -6350 15350
rect -6300 15300 -5800 18700
rect -9700 14800 -5800 15300
rect -6300 14750 -5800 14800
rect -5750 14750 -5250 18700
rect -9700 14250 -5250 14750
rect -5750 14200 -5250 14250
rect -5200 14200 -4700 18700
rect -9700 13700 -4700 14200
rect -5200 13650 -4700 13700
rect -4650 13650 -4150 18700
rect -9700 13150 -4150 13650
rect -4650 13100 -4150 13150
rect -4100 13100 -3600 18700
rect -9700 12600 -3600 13100
rect -4100 12550 -3600 12600
rect -3550 12550 -3050 18700
rect -9700 12050 -3050 12550
rect -3550 12000 -3050 12050
rect -3000 12000 -2500 18700
rect -9700 11500 -2500 12000
rect -3000 11450 -2500 11500
rect -2450 11450 -1950 18700
rect -9700 10950 -1950 11450
rect -2450 10900 -1950 10950
rect -1900 10900 -1400 18700
rect -9700 10400 -1400 10900
rect -1900 10350 -1400 10400
rect -1350 10350 -850 18700
rect -9700 9850 -850 10350
rect -1350 9800 -850 9850
rect -800 9800 -300 18700
rect -9700 9300 -300 9800
rect -800 9250 -300 9300
rect -250 9250 250 18700
rect 300 9800 800 18700
rect 850 10350 1350 18700
rect 1400 10900 1900 18700
rect 1950 11450 2450 18700
rect 2500 12000 3000 18700
rect 3050 12550 3550 18700
rect 3600 13100 4100 18700
rect 4150 13650 4650 18700
rect 4700 14200 5200 18700
rect 5250 14750 5750 18700
rect 5800 15300 6300 18700
rect 6350 15850 6850 18700
rect 6900 16400 7400 18700
rect 7450 16950 7950 18700
rect 8000 17500 8500 18700
rect 8000 17000 9700 17500
rect 8000 16950 8500 17000
rect 7450 16450 9700 16950
rect 7450 16400 7950 16450
rect 6900 15900 9700 16400
rect 6900 15850 7400 15900
rect 6350 15350 9700 15850
rect 6350 15300 6850 15350
rect 5800 14800 9700 15300
rect 5800 14750 6300 14800
rect 5250 14250 9700 14750
rect 5250 14200 5750 14250
rect 4700 13700 9700 14200
rect 4700 13650 5200 13700
rect 4150 13150 9700 13650
rect 4150 13100 4650 13150
rect 3600 12600 9700 13100
rect 3600 12550 4100 12600
rect 3050 12050 9700 12550
rect 3050 12000 3550 12050
rect 2500 11500 9700 12000
rect 2500 11450 3000 11500
rect 1950 10950 9700 11450
rect 1950 10900 2450 10950
rect 1400 10400 9700 10900
rect 1400 10350 1900 10400
rect 850 9850 9700 10350
rect 850 9800 1350 9850
rect 300 9300 9700 9800
rect 300 9250 800 9300
rect -9700 9230 9700 9250
rect -9700 8750 -230 9230
rect -250 8700 -230 8750
rect -9750 8200 -230 8700
rect -250 8150 -230 8200
rect -9700 7670 -230 8150
rect 230 8750 9700 9230
rect 230 8700 250 8750
rect 230 8200 9700 8700
rect 230 8150 250 8200
rect 230 7670 9700 8150
rect -9700 7650 9700 7670
rect -800 7600 -300 7650
rect -9700 7100 -300 7600
rect -1350 7050 -850 7100
rect -9700 6550 -850 7050
rect -1900 6500 -1400 6550
rect -9700 6000 -1400 6500
rect -2450 5950 -1950 6000
rect -9700 5450 -1950 5950
rect -3000 5400 -2500 5450
rect -9700 4900 -2500 5400
rect -3550 4850 -3050 4900
rect -9700 4350 -3050 4850
rect -4100 4300 -3600 4350
rect -9700 3800 -3600 4300
rect -4650 3750 -4150 3800
rect -9700 3250 -4150 3750
rect -5200 3200 -4700 3250
rect -9700 2700 -4700 3200
rect -5750 2650 -5250 2700
rect -9700 2150 -5250 2650
rect -6300 2100 -5800 2150
rect -9700 1600 -5800 2100
rect -6850 1550 -6350 1600
rect -9700 1050 -6350 1550
rect -7400 1000 -6900 1050
rect -9700 500 -6900 1000
rect -7950 450 -7450 500
rect -9700 -50 -7450 450
rect -8500 -1200 -8000 -50
rect -7950 -1200 -7450 -50
rect -7400 -1200 -6900 500
rect -6850 -1200 -6350 1050
rect -6300 -1200 -5800 1600
rect -5750 -1200 -5250 2150
rect -5200 -1200 -4700 2700
rect -4650 -1200 -4150 3250
rect -4100 -1200 -3600 3800
rect -3550 -1200 -3050 4350
rect -3000 -1200 -2500 4900
rect -2450 -1200 -1950 5450
rect -1900 -1200 -1400 6000
rect -1350 -1200 -850 6550
rect -800 -1200 -300 7100
rect -250 -1200 250 7650
rect 300 7600 800 7650
rect 300 7100 9700 7600
rect 300 -1200 800 7100
rect 850 7050 1350 7100
rect 850 6550 9700 7050
rect 850 -1200 1350 6550
rect 1400 6500 1900 6550
rect 1400 6000 9700 6500
rect 1400 -1200 1900 6000
rect 1950 5950 2450 6000
rect 1950 5450 9700 5950
rect 1950 -1200 2450 5450
rect 2500 5400 3000 5450
rect 2500 4900 9700 5400
rect 2500 -1200 3000 4900
rect 3050 4850 3550 4900
rect 3050 4350 9700 4850
rect 3050 -1200 3550 4350
rect 3600 4300 4100 4350
rect 3600 3800 9700 4300
rect 3600 -1200 4100 3800
rect 4150 3750 4650 3800
rect 4150 3250 9700 3750
rect 4150 -1200 4650 3250
rect 4700 3200 5200 3250
rect 4700 2700 9700 3200
rect 4700 -1200 5200 2700
rect 5250 2650 5750 2700
rect 5250 2150 9700 2650
rect 5250 -1200 5750 2150
rect 5800 2100 6300 2150
rect 5800 1600 9700 2100
rect 5800 -1200 6300 1600
rect 6350 1550 6850 1600
rect 6350 1050 9700 1550
rect 6350 -1200 6850 1050
rect 6900 1000 7400 1050
rect 6900 500 9700 1000
rect 6900 -1200 7400 500
rect 7450 450 7950 500
rect 7450 -50 9700 450
rect 7450 -1200 7950 -50
rect 8000 -1200 8500 -50
<< viali >>
rect -230 7670 230 9230
<< metal1 >>
rect -250 9230 250 9250
rect -250 7670 -230 9230
rect 230 7670 250 9230
rect -250 -1500 250 7670
<< metal4 >>
rect -3728 18400 -493 18500
rect -3728 17600 -3628 18400
rect -1300 18000 -493 18400
tri -493 18000 7 18500 sw
rect -1300 17600 7 18000
rect -3728 17500 7 17600
tri -907 16586 7 17500 ne
tri 7 17100 907 18000 sw
rect 7 17000 3148 17100
rect 7 16586 1300 17000
tri 7 16100 493 16586 ne
rect 493 16200 1300 16586
rect 3048 16200 3148 17000
rect 493 16100 3148 16200
<< via4 >>
rect -3628 17600 -1300 18400
rect 1300 16200 3048 17000
<< metal5 >>
tri -5335 17100 -3935 18500 se
rect -3935 18400 -1200 18500
rect -3935 17600 -3628 18400
rect -1300 17600 -1200 18400
rect -3935 17500 -1200 17600
rect -3935 17100 -3921 17500
tri -3921 17100 -3521 17500 nw
tri -907 17100 493 18500 se
rect 493 18000 3935 18500
tri 3935 18000 4435 18500 sw
rect 493 17500 4435 18000
rect 493 17100 507 17500
tri 507 17100 907 17500 nw
tri 3521 17100 3921 17500 ne
rect 3921 17100 4435 17500
tri -6556 15879 -5335 17100 se
rect -5335 16727 -4294 17100
tri -4294 16727 -3921 17100 nw
tri -3728 16727 -3355 17100 se
rect -3355 16727 -493 17100
rect -5335 16459 -4562 16727
tri -4562 16459 -4294 16727 nw
tri -3996 16459 -3728 16727 se
rect -3728 16459 -493 16727
rect -5335 15893 -5128 16459
tri -5128 15893 -4562 16459 nw
tri -4562 15893 -3996 16459 se
rect -3996 16100 -493 16459
tri -493 16100 507 17100 nw
rect 1200 17000 3355 17100
rect 1200 16200 1300 17000
rect 3048 16586 3355 17000
tri 3355 16586 3869 17100 sw
tri 3921 16586 4435 17100 ne
tri 4435 16586 5849 18000 sw
rect 3048 16200 3869 16586
rect 1200 16100 3869 16200
rect -3996 15893 -3162 16100
rect -5335 15879 -5142 15893
tri -5142 15879 -5128 15893 nw
tri -4576 15879 -4562 15893 se
rect -4562 15879 -3162 15893
tri -3162 15879 -2941 16100 nw
tri -7970 14465 -6556 15879 se
rect -6556 15313 -5708 15879
tri -5708 15313 -5142 15879 nw
tri -5142 15313 -4576 15879 se
rect -6556 15045 -5976 15313
tri -5976 15045 -5708 15313 nw
tri -5410 15045 -5142 15313 se
rect -5142 15045 -4576 15313
rect -6556 14479 -6542 15045
tri -6542 14479 -5976 15045 nw
tri -5976 14479 -5410 15045 se
rect -5410 14479 -4576 15045
tri -6556 14465 -6542 14479 nw
tri -5990 14465 -5976 14479 se
rect -5976 14465 -4576 14479
tri -4576 14465 -3162 15879 nw
tri 2941 15172 3869 16100 ne
tri 3869 16020 4435 16586 sw
tri 4435 16020 5001 16586 ne
rect 5001 16020 5849 16586
rect 3869 15752 4435 16020
tri 4435 15752 4703 16020 sw
tri 5001 15752 5269 16020 ne
rect 5269 15752 5849 16020
rect 3869 15186 4703 15752
tri 4703 15186 5269 15752 sw
tri 5269 15186 5835 15752 ne
rect 5835 15186 5849 15752
rect 3869 15172 5269 15186
tri 5269 15172 5283 15186 sw
tri 5835 15172 5849 15186 ne
tri 5849 15172 7263 16586 sw
tri -9384 13051 -7970 14465 se
rect -7970 13899 -7122 14465
tri -7122 13899 -6556 14465 nw
tri -6556 13899 -5990 14465 se
rect -7970 13631 -7390 13899
tri -7390 13631 -7122 13899 nw
tri -6824 13631 -6556 13899 se
rect -6556 13631 -5990 13899
rect -7970 13065 -7956 13631
tri -7956 13065 -7390 13631 nw
tri -7390 13065 -6824 13631 se
rect -6824 13065 -5990 13631
tri -7970 13051 -7956 13065 nw
tri -7404 13051 -7390 13065 se
rect -7390 13051 -5990 13065
tri -5990 13051 -4576 14465 nw
tri 3869 13758 5283 15172 ne
tri 5283 14606 5849 15172 sw
tri 5849 14606 6415 15172 ne
rect 6415 14606 7263 15172
rect 5283 14338 5849 14606
tri 5849 14338 6117 14606 sw
tri 6415 14338 6683 14606 ne
rect 6683 14338 7263 14606
rect 5283 13772 6117 14338
tri 6117 13772 6683 14338 sw
tri 6683 13772 7249 14338 ne
rect 7249 13772 7263 14338
rect 5283 13758 6683 13772
tri 6683 13758 6697 13772 sw
tri 7249 13758 7263 13772 ne
tri 7263 13758 8677 15172 sw
tri -9500 12935 -9384 13051 se
rect -9384 12935 -8500 13051
rect -9500 5105 -8500 12935
tri -8500 12521 -7970 13051 nw
tri -7970 12485 -7404 13051 se
rect -7404 12485 -7100 13051
tri -8100 12355 -7970 12485 se
rect -7970 12355 -7100 12485
rect -8100 5645 -7100 12355
tri -7100 11941 -5990 13051 nw
tri 5283 12358 6683 13758 ne
rect 6683 13192 6697 13758
tri 6697 13192 7263 13758 sw
tri 7263 13192 7829 13758 ne
rect 7829 13192 8677 13758
rect 6683 12924 7263 13192
tri 7263 12924 7531 13192 sw
tri 7829 12924 8097 13192 ne
rect 8097 12935 8677 13192
tri 8677 12935 9500 13758 sw
rect 8097 12924 9500 12935
rect 6683 12358 7531 12924
tri 7531 12358 8097 12924 sw
tri 8097 12521 8500 12924 ne
tri 6683 11941 7100 12358 ne
rect 7100 12355 8097 12358
tri 8097 12355 8100 12358 sw
tri -8500 5105 -8126 5479 sw
tri -8100 5105 -7560 5645 ne
rect -7560 5642 -7100 5645
tri -7100 5642 -6683 6059 sw
tri 6893 5852 7100 6059 se
rect 7100 5852 8100 12355
rect -7560 5105 -6683 5642
rect -9500 5065 -8126 5105
tri -9500 4242 -8677 5065 ne
rect -8677 4808 -8126 5065
tri -8126 4808 -7829 5105 sw
tri -7560 4808 -7263 5105 ne
rect -7263 4808 -6683 5105
rect -8677 4242 -7829 4808
tri -7829 4242 -7263 4808 sw
tri -7263 4242 -6697 4808 ne
rect -6697 4242 -6683 4808
tri -8677 2828 -7263 4242 ne
tri -7263 4228 -7249 4242 sw
tri -6697 4228 -6683 4242 ne
tri -6683 4228 -5269 5642 sw
tri 5976 4935 6893 5852 se
rect 6893 5645 8100 5852
rect 6893 5272 7727 5645
tri 7727 5272 8100 5645 nw
tri 8293 5272 8500 5479 se
rect 8500 5272 9500 12924
rect 6893 4935 7390 5272
tri 7390 4935 7727 5272 nw
tri 7956 4935 8293 5272 se
rect 8293 5065 9500 5272
rect 8293 4935 9370 5065
tri 9370 4935 9500 5065 nw
rect -7263 3662 -7249 4228
tri -7249 3662 -6683 4228 sw
tri -6683 3662 -6117 4228 ne
rect -6117 3662 -5269 4228
rect -7263 3394 -6683 3662
tri -6683 3394 -6415 3662 sw
tri -6117 3394 -5849 3662 ne
rect -5849 3394 -5269 3662
rect -7263 2828 -6415 3394
tri -6415 2828 -5849 3394 sw
tri -5849 2828 -5283 3394 ne
rect -5283 2828 -5269 3394
tri -7263 1414 -5849 2828 ne
tri -5849 2814 -5835 2828 sw
tri -5283 2814 -5269 2828 ne
tri -5269 2814 -3855 4228 sw
tri 4562 3521 5976 4935 se
rect 5976 4369 6824 4935
tri 6824 4369 7390 4935 nw
tri 7390 4369 7956 4935 se
rect 5976 4101 6556 4369
tri 6556 4101 6824 4369 nw
tri 7122 4101 7390 4369 se
rect 7390 4101 7956 4369
rect 5976 3535 5990 4101
tri 5990 3535 6556 4101 nw
tri 6556 3535 7122 4101 se
rect 7122 3535 7956 4101
tri 5976 3521 5990 3535 nw
tri 6542 3521 6556 3535 se
rect 6556 3521 7956 3535
tri 7956 3521 9370 4935 nw
rect -5849 2248 -5835 2814
tri -5835 2248 -5269 2814 sw
tri -5269 2248 -4703 2814 ne
rect -4703 2248 -3855 2814
rect -5849 1980 -5269 2248
tri -5269 1980 -5001 2248 sw
tri -4703 1980 -4435 2248 ne
rect -4435 1980 -3855 2248
rect -5849 1414 -5001 1980
tri -5001 1414 -4435 1980 sw
tri -4435 1414 -3869 1980 ne
rect -3869 1900 -3855 1980
tri -3855 1900 -2941 2814 sw
tri 3148 2107 4562 3521 se
rect 4562 2955 5410 3521
tri 5410 2955 5976 3521 nw
tri 5976 2955 6542 3521 se
rect 4562 2687 5142 2955
tri 5142 2687 5410 2955 nw
tri 5708 2687 5976 2955 se
rect 5976 2687 6542 2955
rect 4562 2121 4576 2687
tri 4576 2121 5142 2687 nw
tri 5142 2121 5708 2687 se
rect 5708 2121 6542 2687
tri 4562 2107 4576 2121 nw
tri 5128 2107 5142 2121 se
rect 5142 2107 6542 2121
tri 6542 2107 7956 3521 nw
tri 2941 1900 3148 2107 se
rect 3148 1900 3996 2107
rect -3869 1541 3996 1900
tri 3996 1541 4562 2107 nw
tri 4562 1541 5128 2107 se
rect 5128 1541 5142 2107
rect -3869 1414 3728 1541
tri -5849 0 -4435 1414 ne
tri -4435 900 -3921 1414 sw
tri -3869 900 -3355 1414 ne
rect -3355 1273 3728 1414
tri 3728 1273 3996 1541 nw
tri 4294 1273 4562 1541 se
rect 4562 1273 5142 1541
rect -3355 900 3355 1273
tri 3355 900 3728 1273 nw
rect -4435 500 -3921 900
tri -3921 500 -3521 900 sw
rect -4435 0 -2728 500
tri -4435 -500 -3935 0 ne
rect -3935 -500 -2728 0
rect -3728 -1500 -2728 -500
rect -500 -1500 500 900
tri 3728 707 4294 1273 se
rect 4294 707 5142 1273
tri 5142 707 6542 2107 nw
tri 3521 500 3728 707 se
rect 3728 500 3935 707
rect 2728 -500 3935 500
tri 3935 -500 5142 707 nw
rect 2728 -1500 3728 -500
<< end >>
