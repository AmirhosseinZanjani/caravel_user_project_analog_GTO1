magic
tech sky130A
magscale 1 2
timestamp 1695391617
<< pwell >>
rect -134 188 -24 938
rect 1050 188 1160 938
rect 30 14 96 150
rect 921 109 927 161
rect 930 14 996 150
<< locali >>
rect -134 188 16 938
rect 1010 188 1160 938
rect 30 14 96 150
rect 930 14 996 150
<< metal1 >>
rect -87 1444 -39 1562
rect -89 1438 -37 1444
rect -89 1380 -37 1386
rect -87 -62 -39 1380
rect 9 1252 57 1562
rect 105 1540 153 1562
rect 103 1534 155 1540
rect 103 1476 155 1482
rect 7 1246 59 1252
rect 7 1188 59 1194
rect 9 926 57 1188
rect 105 926 153 1476
rect 201 1348 249 1562
rect 199 1342 251 1348
rect 199 1284 251 1290
rect 201 926 249 1284
rect 297 1252 345 1562
rect 393 1348 441 1562
rect 489 1540 537 1562
rect 487 1534 539 1540
rect 487 1476 539 1482
rect 489 1444 537 1476
rect 487 1438 539 1444
rect 487 1380 539 1386
rect 391 1342 443 1348
rect 391 1284 443 1290
rect 295 1246 347 1252
rect 295 1188 347 1194
rect 297 926 345 1188
rect 393 926 441 1284
rect 489 926 537 1380
rect 585 1348 633 1562
rect 583 1342 635 1348
rect 583 1284 635 1290
rect 585 926 633 1284
rect 681 1252 729 1562
rect 777 1348 825 1562
rect 873 1444 921 1562
rect 871 1438 923 1444
rect 871 1380 923 1386
rect 775 1342 827 1348
rect 775 1284 827 1290
rect 679 1246 731 1252
rect 679 1188 731 1194
rect 681 926 729 1188
rect 777 926 825 1284
rect 873 926 921 1380
rect 969 1252 1017 1562
rect 1065 1540 1113 1562
rect 1063 1534 1115 1540
rect 1063 1476 1115 1482
rect 967 1246 1019 1252
rect 967 1188 1019 1194
rect 969 926 1017 1188
rect 105 110 206 156
rect 258 110 345 156
rect 369 110 384 156
rect 450 110 576 156
rect 642 110 768 156
rect 820 110 921 156
rect 105 -62 153 110
rect -89 -68 -37 -62
rect -89 -126 -37 -120
rect 103 -68 155 -62
rect 103 -126 155 -120
rect -87 -225 -39 -126
rect 105 -225 153 -126
rect 297 -158 345 110
rect 489 -62 537 110
rect 487 -68 539 -62
rect 487 -126 539 -120
rect 295 -164 347 -158
rect 295 -222 347 -216
rect 297 -225 345 -222
rect 489 -225 537 -126
rect 681 -158 729 110
rect 873 -62 921 110
rect 1065 -62 1113 1476
rect 871 -68 923 -62
rect 871 -126 923 -120
rect 1063 -68 1115 -62
rect 1063 -126 1115 -120
rect 679 -164 731 -158
rect 679 -222 731 -216
rect 681 -225 729 -222
rect 873 -225 921 -126
rect 1065 -225 1113 -126
<< via1 >>
rect -89 1386 -37 1438
rect 103 1482 155 1534
rect 7 1194 59 1246
rect 199 1290 251 1342
rect 487 1482 539 1534
rect 487 1386 539 1438
rect 391 1290 443 1342
rect 295 1194 347 1246
rect 583 1290 635 1342
rect 871 1386 923 1438
rect 775 1290 827 1342
rect 679 1194 731 1246
rect 1063 1482 1115 1534
rect 967 1194 1019 1246
rect -89 -120 -37 -68
rect 103 -120 155 -68
rect 487 -120 539 -68
rect 295 -216 347 -164
rect 871 -120 923 -68
rect 1063 -120 1115 -68
rect 679 -216 731 -164
<< metal2 >>
rect 103 1534 155 1540
rect -134 1484 103 1532
rect 487 1534 539 1540
rect 155 1484 487 1532
rect 103 1476 155 1482
rect 487 1476 539 1482
rect 1063 1534 1115 1540
rect 1115 1484 1160 1532
rect 1063 1476 1115 1482
rect -89 1438 -37 1444
rect -134 1388 -89 1436
rect -89 1380 -37 1386
rect 487 1438 539 1444
rect 871 1438 923 1444
rect 539 1388 871 1436
rect 487 1380 539 1386
rect 923 1388 1160 1436
rect 871 1380 923 1386
rect 199 1342 251 1348
rect -94 1292 199 1340
rect 391 1342 443 1348
rect 251 1292 391 1340
rect 199 1284 251 1290
rect 583 1342 635 1348
rect 443 1292 583 1340
rect 391 1284 443 1290
rect 775 1342 827 1348
rect 635 1292 775 1340
rect 583 1284 635 1290
rect 827 1292 1118 1340
rect 775 1284 827 1290
rect 7 1246 59 1252
rect -94 1196 7 1244
rect 295 1246 347 1252
rect 59 1196 295 1244
rect 7 1188 59 1194
rect 679 1246 731 1252
rect 347 1196 679 1244
rect 295 1188 347 1194
rect 967 1246 1019 1252
rect 731 1196 967 1244
rect 679 1188 731 1194
rect 1019 1196 1118 1244
rect 967 1188 1019 1194
rect -89 -68 -37 -62
rect -94 -118 -89 -70
rect 103 -68 155 -62
rect -37 -118 103 -70
rect -89 -126 -37 -120
rect 487 -68 539 -62
rect 155 -118 487 -70
rect 103 -126 155 -120
rect 871 -68 923 -62
rect 539 -118 871 -70
rect 487 -126 539 -120
rect 1063 -68 1115 -62
rect 923 -118 1063 -70
rect 871 -126 923 -120
rect 1115 -118 1120 -70
rect 1063 -126 1115 -120
rect 295 -164 347 -158
rect -134 -214 295 -166
rect 679 -164 731 -158
rect 347 -214 679 -166
rect 295 -222 347 -216
rect 731 -214 1160 -166
rect 679 -222 731 -216
use sky130_fd_pr__nfet_01v8_QMBXET  sky130_fd_pr__nfet_01v8_QMBXET_0
timestamp 1695389752
transform 1 0 513 0 1 563
box -647 -585 647 585
<< labels >>
flabel locali -134 188 16 938 0 FreeSans 320 0 0 0 VSUB
port 0 nsew
flabel locali 1010 188 1160 938 0 FreeSans 320 0 0 0 VSUB
port 0 nsew
flabel metal2 -134 1484 -89 1532 0 FreeSans 128 0 0 0 drain
port 2 nsew
flabel metal2 -134 -214 -88 -166 0 FreeSans 128 0 0 0 en
port 3 nsew
flabel metal2 -134 1388 -89 1436 0 FreeSans 128 0 0 0 gate
port 1 nsew
<< end >>
