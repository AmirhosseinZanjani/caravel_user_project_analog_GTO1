magic
tech sky130A
magscale 1 2
timestamp 1695283740
<< error_s >>
rect 47 137 105 143
rect 1331 137 1389 143
rect 47 103 59 137
rect 1331 103 1343 137
rect 47 97 105 103
rect 1331 97 1389 103
<< locali >>
rect 1370 184 1522 666
rect 48 3 104 137
rect 1332 3 1388 137
<< metal1 >>
rect 118 1182 166 1190
rect 116 1176 168 1182
rect 116 1118 168 1124
rect 118 674 166 1118
rect 214 1086 262 1190
rect 212 1080 264 1086
rect 212 1022 264 1028
rect 214 674 262 1022
rect 310 990 358 1190
rect 406 1086 454 1190
rect 502 1182 550 1190
rect 500 1176 552 1182
rect 500 1118 552 1124
rect 404 1080 456 1086
rect 404 1022 456 1028
rect 308 984 360 990
rect 308 926 360 932
rect 310 674 358 926
rect 406 674 454 1022
rect 502 674 550 1118
rect 598 1086 646 1190
rect 596 1080 648 1086
rect 596 1022 648 1028
rect 598 674 646 1022
rect 694 990 742 1190
rect 790 1086 838 1190
rect 886 1182 934 1190
rect 884 1176 936 1182
rect 884 1118 936 1124
rect 788 1080 840 1086
rect 788 1022 840 1028
rect 692 984 744 990
rect 692 926 744 932
rect 694 674 742 926
rect 790 674 838 1022
rect 886 674 934 1118
rect 982 1086 1030 1190
rect 980 1080 1032 1086
rect 980 1022 1032 1028
rect 982 674 1030 1022
rect 1078 990 1126 1190
rect 1174 1086 1222 1190
rect 1270 1182 1318 1190
rect 1268 1176 1320 1182
rect 1268 1118 1320 1124
rect 1172 1080 1224 1086
rect 1172 1022 1224 1028
rect 1076 984 1128 990
rect 1076 926 1128 932
rect 1078 674 1126 926
rect 1174 674 1222 1022
rect 1270 674 1318 1118
rect 166 -172 214 140
rect 310 -76 358 140
rect 308 -82 360 -76
rect 308 -140 360 -134
rect 164 -178 216 -172
rect 164 -236 216 -230
rect 166 -246 214 -236
rect 310 -244 358 -140
rect 502 -172 550 140
rect 694 -76 742 140
rect 692 -82 744 -76
rect 692 -140 744 -134
rect 500 -178 552 -172
rect 500 -236 552 -230
rect 502 -246 550 -236
rect 694 -244 742 -140
rect 886 -172 934 140
rect 1078 -76 1126 140
rect 1076 -82 1128 -76
rect 1076 -140 1128 -134
rect 884 -178 936 -172
rect 884 -236 936 -230
rect 886 -244 934 -236
rect 1078 -244 1126 -140
rect 1222 -172 1270 140
rect 1220 -178 1272 -172
rect 1220 -236 1272 -230
rect 1222 -244 1270 -236
<< via1 >>
rect 116 1124 168 1176
rect 212 1028 264 1080
rect 500 1124 552 1176
rect 404 1028 456 1080
rect 308 932 360 984
rect 596 1028 648 1080
rect 884 1124 936 1176
rect 788 1028 840 1080
rect 692 932 744 984
rect 980 1028 1032 1080
rect 1268 1124 1320 1176
rect 1172 1028 1224 1080
rect 1076 932 1128 984
rect 308 -134 360 -82
rect 164 -230 216 -178
rect 692 -134 744 -82
rect 500 -230 552 -178
rect 1076 -134 1128 -82
rect 884 -230 936 -178
rect 1220 -230 1272 -178
<< metal2 >>
rect 116 1176 168 1182
rect -122 1126 116 1174
rect 500 1176 552 1182
rect 168 1126 500 1174
rect 116 1118 168 1124
rect 884 1176 936 1182
rect 552 1126 884 1174
rect 500 1118 552 1124
rect 1268 1176 1320 1182
rect 936 1126 1268 1174
rect 884 1118 936 1124
rect 1320 1126 1558 1174
rect 1268 1118 1320 1124
rect 212 1080 264 1086
rect -122 1030 212 1078
rect 404 1080 456 1086
rect 264 1030 404 1078
rect 212 1022 264 1028
rect 596 1080 648 1086
rect 456 1030 596 1078
rect 404 1022 456 1028
rect 788 1080 840 1086
rect 648 1030 788 1078
rect 596 1022 648 1028
rect 980 1080 1032 1086
rect 840 1030 980 1078
rect 788 1022 840 1028
rect 1172 1080 1224 1086
rect 1032 1030 1172 1078
rect 980 1022 1032 1028
rect 1224 1030 1558 1078
rect 1172 1022 1224 1028
rect 308 984 360 990
rect -122 934 308 982
rect 692 984 744 990
rect 360 934 692 982
rect 308 926 360 932
rect 1076 984 1128 990
rect 744 934 1076 982
rect 692 926 744 932
rect 1128 934 1558 982
rect 1076 926 1128 932
rect 308 -82 360 -76
rect -122 -132 308 -84
rect 692 -82 744 -76
rect 360 -132 692 -84
rect 308 -140 360 -134
rect 1076 -82 1128 -76
rect 744 -132 1076 -84
rect 692 -140 744 -134
rect 1128 -132 1558 -84
rect 1076 -140 1128 -134
rect 164 -178 216 -172
rect -122 -228 164 -180
rect 500 -178 552 -172
rect 216 -228 500 -180
rect 164 -236 216 -230
rect 884 -178 936 -172
rect 552 -228 884 -180
rect 500 -236 552 -230
rect 1220 -178 1272 -172
rect 936 -228 1220 -180
rect 884 -236 936 -230
rect 1272 -228 1558 -180
rect 1220 -236 1272 -230
use sky130_fd_pr__nfet_01v8_LM9D52  sky130_fd_pr__nfet_01v8_LM9D52_0
timestamp 1694525365
transform 1 0 718 0 1 425
box -839 -460 839 460
<< labels >>
flabel metal2 -122 1030 116 1078 0 FreeSans 320 0 160 0 M1S_M2D
flabel metal2 -122 1126 1558 1174 0 FreeSans 320 0 -6240 0 M2S
flabel metal2 -122 934 692 982 0 FreeSans 320 0 -2720 0 M1D
flabel metal2 -122 -132 308 -84 0 FreeSans 320 0 -1120 0 M1G
flabel metal2 -122 -228 164 -180 0 FreeSans 320 0 -480 0 M2G
rlabel metal2 -122 -204 -122 -204 3 M2G
port 2 e
rlabel metal2 -122 -108 -122 -108 3 M1G
port 1 e
rlabel metal2 -122 958 -122 958 3 M1D
port 3 e
rlabel metal2 -122 1056 -122 1056 3 M1S_M2D
port 4 e
rlabel metal2 -122 1150 -122 1150 3 M2S
port 5 e
<< end >>
