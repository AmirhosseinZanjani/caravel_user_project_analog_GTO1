magic
tech sky130A
magscale 1 2
timestamp 1693317617
<< pwell >>
rect -4037 -310 4037 310
<< nmos >>
rect -3841 -100 -3641 100
rect -3583 -100 -3383 100
rect -3325 -100 -3125 100
rect -3067 -100 -2867 100
rect -2809 -100 -2609 100
rect -2551 -100 -2351 100
rect -2293 -100 -2093 100
rect -2035 -100 -1835 100
rect -1777 -100 -1577 100
rect -1519 -100 -1319 100
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
rect 1319 -100 1519 100
rect 1577 -100 1777 100
rect 1835 -100 2035 100
rect 2093 -100 2293 100
rect 2351 -100 2551 100
rect 2609 -100 2809 100
rect 2867 -100 3067 100
rect 3125 -100 3325 100
rect 3383 -100 3583 100
rect 3641 -100 3841 100
<< ndiff >>
rect -3899 88 -3841 100
rect -3899 -88 -3887 88
rect -3853 -88 -3841 88
rect -3899 -100 -3841 -88
rect -3641 88 -3583 100
rect -3641 -88 -3629 88
rect -3595 -88 -3583 88
rect -3641 -100 -3583 -88
rect -3383 88 -3325 100
rect -3383 -88 -3371 88
rect -3337 -88 -3325 88
rect -3383 -100 -3325 -88
rect -3125 88 -3067 100
rect -3125 -88 -3113 88
rect -3079 -88 -3067 88
rect -3125 -100 -3067 -88
rect -2867 88 -2809 100
rect -2867 -88 -2855 88
rect -2821 -88 -2809 88
rect -2867 -100 -2809 -88
rect -2609 88 -2551 100
rect -2609 -88 -2597 88
rect -2563 -88 -2551 88
rect -2609 -100 -2551 -88
rect -2351 88 -2293 100
rect -2351 -88 -2339 88
rect -2305 -88 -2293 88
rect -2351 -100 -2293 -88
rect -2093 88 -2035 100
rect -2093 -88 -2081 88
rect -2047 -88 -2035 88
rect -2093 -100 -2035 -88
rect -1835 88 -1777 100
rect -1835 -88 -1823 88
rect -1789 -88 -1777 88
rect -1835 -100 -1777 -88
rect -1577 88 -1519 100
rect -1577 -88 -1565 88
rect -1531 -88 -1519 88
rect -1577 -100 -1519 -88
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
rect 1519 88 1577 100
rect 1519 -88 1531 88
rect 1565 -88 1577 88
rect 1519 -100 1577 -88
rect 1777 88 1835 100
rect 1777 -88 1789 88
rect 1823 -88 1835 88
rect 1777 -100 1835 -88
rect 2035 88 2093 100
rect 2035 -88 2047 88
rect 2081 -88 2093 88
rect 2035 -100 2093 -88
rect 2293 88 2351 100
rect 2293 -88 2305 88
rect 2339 -88 2351 88
rect 2293 -100 2351 -88
rect 2551 88 2609 100
rect 2551 -88 2563 88
rect 2597 -88 2609 88
rect 2551 -100 2609 -88
rect 2809 88 2867 100
rect 2809 -88 2821 88
rect 2855 -88 2867 88
rect 2809 -100 2867 -88
rect 3067 88 3125 100
rect 3067 -88 3079 88
rect 3113 -88 3125 88
rect 3067 -100 3125 -88
rect 3325 88 3383 100
rect 3325 -88 3337 88
rect 3371 -88 3383 88
rect 3325 -100 3383 -88
rect 3583 88 3641 100
rect 3583 -88 3595 88
rect 3629 -88 3641 88
rect 3583 -100 3641 -88
rect 3841 88 3899 100
rect 3841 -88 3853 88
rect 3887 -88 3899 88
rect 3841 -100 3899 -88
<< ndiffc >>
rect -3887 -88 -3853 88
rect -3629 -88 -3595 88
rect -3371 -88 -3337 88
rect -3113 -88 -3079 88
rect -2855 -88 -2821 88
rect -2597 -88 -2563 88
rect -2339 -88 -2305 88
rect -2081 -88 -2047 88
rect -1823 -88 -1789 88
rect -1565 -88 -1531 88
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect 1531 -88 1565 88
rect 1789 -88 1823 88
rect 2047 -88 2081 88
rect 2305 -88 2339 88
rect 2563 -88 2597 88
rect 2821 -88 2855 88
rect 3079 -88 3113 88
rect 3337 -88 3371 88
rect 3595 -88 3629 88
rect 3853 -88 3887 88
<< psubdiff >>
rect -4001 240 -3905 274
rect 3905 240 4001 274
rect -4001 178 -3967 240
rect 3967 178 4001 240
rect -4001 -240 -3967 -178
rect 3967 -240 4001 -178
rect -4001 -274 -3905 -240
rect 3905 -274 4001 -240
<< psubdiffcont >>
rect -3905 240 3905 274
rect -4001 -178 -3967 178
rect 3967 -178 4001 178
rect -3905 -274 3905 -240
<< poly >>
rect -3841 172 -3641 188
rect -3841 138 -3825 172
rect -3657 138 -3641 172
rect -3841 100 -3641 138
rect -3583 172 -3383 188
rect -3583 138 -3567 172
rect -3399 138 -3383 172
rect -3583 100 -3383 138
rect -3325 172 -3125 188
rect -3325 138 -3309 172
rect -3141 138 -3125 172
rect -3325 100 -3125 138
rect -3067 172 -2867 188
rect -3067 138 -3051 172
rect -2883 138 -2867 172
rect -3067 100 -2867 138
rect -2809 172 -2609 188
rect -2809 138 -2793 172
rect -2625 138 -2609 172
rect -2809 100 -2609 138
rect -2551 172 -2351 188
rect -2551 138 -2535 172
rect -2367 138 -2351 172
rect -2551 100 -2351 138
rect -2293 172 -2093 188
rect -2293 138 -2277 172
rect -2109 138 -2093 172
rect -2293 100 -2093 138
rect -2035 172 -1835 188
rect -2035 138 -2019 172
rect -1851 138 -1835 172
rect -2035 100 -1835 138
rect -1777 172 -1577 188
rect -1777 138 -1761 172
rect -1593 138 -1577 172
rect -1777 100 -1577 138
rect -1519 172 -1319 188
rect -1519 138 -1503 172
rect -1335 138 -1319 172
rect -1519 100 -1319 138
rect -1261 172 -1061 188
rect -1261 138 -1245 172
rect -1077 138 -1061 172
rect -1261 100 -1061 138
rect -1003 172 -803 188
rect -1003 138 -987 172
rect -819 138 -803 172
rect -1003 100 -803 138
rect -745 172 -545 188
rect -745 138 -729 172
rect -561 138 -545 172
rect -745 100 -545 138
rect -487 172 -287 188
rect -487 138 -471 172
rect -303 138 -287 172
rect -487 100 -287 138
rect -229 172 -29 188
rect -229 138 -213 172
rect -45 138 -29 172
rect -229 100 -29 138
rect 29 172 229 188
rect 29 138 45 172
rect 213 138 229 172
rect 29 100 229 138
rect 287 172 487 188
rect 287 138 303 172
rect 471 138 487 172
rect 287 100 487 138
rect 545 172 745 188
rect 545 138 561 172
rect 729 138 745 172
rect 545 100 745 138
rect 803 172 1003 188
rect 803 138 819 172
rect 987 138 1003 172
rect 803 100 1003 138
rect 1061 172 1261 188
rect 1061 138 1077 172
rect 1245 138 1261 172
rect 1061 100 1261 138
rect 1319 172 1519 188
rect 1319 138 1335 172
rect 1503 138 1519 172
rect 1319 100 1519 138
rect 1577 172 1777 188
rect 1577 138 1593 172
rect 1761 138 1777 172
rect 1577 100 1777 138
rect 1835 172 2035 188
rect 1835 138 1851 172
rect 2019 138 2035 172
rect 1835 100 2035 138
rect 2093 172 2293 188
rect 2093 138 2109 172
rect 2277 138 2293 172
rect 2093 100 2293 138
rect 2351 172 2551 188
rect 2351 138 2367 172
rect 2535 138 2551 172
rect 2351 100 2551 138
rect 2609 172 2809 188
rect 2609 138 2625 172
rect 2793 138 2809 172
rect 2609 100 2809 138
rect 2867 172 3067 188
rect 2867 138 2883 172
rect 3051 138 3067 172
rect 2867 100 3067 138
rect 3125 172 3325 188
rect 3125 138 3141 172
rect 3309 138 3325 172
rect 3125 100 3325 138
rect 3383 172 3583 188
rect 3383 138 3399 172
rect 3567 138 3583 172
rect 3383 100 3583 138
rect 3641 172 3841 188
rect 3641 138 3657 172
rect 3825 138 3841 172
rect 3641 100 3841 138
rect -3841 -138 -3641 -100
rect -3841 -172 -3825 -138
rect -3657 -172 -3641 -138
rect -3841 -188 -3641 -172
rect -3583 -138 -3383 -100
rect -3583 -172 -3567 -138
rect -3399 -172 -3383 -138
rect -3583 -188 -3383 -172
rect -3325 -138 -3125 -100
rect -3325 -172 -3309 -138
rect -3141 -172 -3125 -138
rect -3325 -188 -3125 -172
rect -3067 -138 -2867 -100
rect -3067 -172 -3051 -138
rect -2883 -172 -2867 -138
rect -3067 -188 -2867 -172
rect -2809 -138 -2609 -100
rect -2809 -172 -2793 -138
rect -2625 -172 -2609 -138
rect -2809 -188 -2609 -172
rect -2551 -138 -2351 -100
rect -2551 -172 -2535 -138
rect -2367 -172 -2351 -138
rect -2551 -188 -2351 -172
rect -2293 -138 -2093 -100
rect -2293 -172 -2277 -138
rect -2109 -172 -2093 -138
rect -2293 -188 -2093 -172
rect -2035 -138 -1835 -100
rect -2035 -172 -2019 -138
rect -1851 -172 -1835 -138
rect -2035 -188 -1835 -172
rect -1777 -138 -1577 -100
rect -1777 -172 -1761 -138
rect -1593 -172 -1577 -138
rect -1777 -188 -1577 -172
rect -1519 -138 -1319 -100
rect -1519 -172 -1503 -138
rect -1335 -172 -1319 -138
rect -1519 -188 -1319 -172
rect -1261 -138 -1061 -100
rect -1261 -172 -1245 -138
rect -1077 -172 -1061 -138
rect -1261 -188 -1061 -172
rect -1003 -138 -803 -100
rect -1003 -172 -987 -138
rect -819 -172 -803 -138
rect -1003 -188 -803 -172
rect -745 -138 -545 -100
rect -745 -172 -729 -138
rect -561 -172 -545 -138
rect -745 -188 -545 -172
rect -487 -138 -287 -100
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -487 -188 -287 -172
rect -229 -138 -29 -100
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect -229 -188 -29 -172
rect 29 -138 229 -100
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 29 -188 229 -172
rect 287 -138 487 -100
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 287 -188 487 -172
rect 545 -138 745 -100
rect 545 -172 561 -138
rect 729 -172 745 -138
rect 545 -188 745 -172
rect 803 -138 1003 -100
rect 803 -172 819 -138
rect 987 -172 1003 -138
rect 803 -188 1003 -172
rect 1061 -138 1261 -100
rect 1061 -172 1077 -138
rect 1245 -172 1261 -138
rect 1061 -188 1261 -172
rect 1319 -138 1519 -100
rect 1319 -172 1335 -138
rect 1503 -172 1519 -138
rect 1319 -188 1519 -172
rect 1577 -138 1777 -100
rect 1577 -172 1593 -138
rect 1761 -172 1777 -138
rect 1577 -188 1777 -172
rect 1835 -138 2035 -100
rect 1835 -172 1851 -138
rect 2019 -172 2035 -138
rect 1835 -188 2035 -172
rect 2093 -138 2293 -100
rect 2093 -172 2109 -138
rect 2277 -172 2293 -138
rect 2093 -188 2293 -172
rect 2351 -138 2551 -100
rect 2351 -172 2367 -138
rect 2535 -172 2551 -138
rect 2351 -188 2551 -172
rect 2609 -138 2809 -100
rect 2609 -172 2625 -138
rect 2793 -172 2809 -138
rect 2609 -188 2809 -172
rect 2867 -138 3067 -100
rect 2867 -172 2883 -138
rect 3051 -172 3067 -138
rect 2867 -188 3067 -172
rect 3125 -138 3325 -100
rect 3125 -172 3141 -138
rect 3309 -172 3325 -138
rect 3125 -188 3325 -172
rect 3383 -138 3583 -100
rect 3383 -172 3399 -138
rect 3567 -172 3583 -138
rect 3383 -188 3583 -172
rect 3641 -138 3841 -100
rect 3641 -172 3657 -138
rect 3825 -172 3841 -138
rect 3641 -188 3841 -172
<< polycont >>
rect -3825 138 -3657 172
rect -3567 138 -3399 172
rect -3309 138 -3141 172
rect -3051 138 -2883 172
rect -2793 138 -2625 172
rect -2535 138 -2367 172
rect -2277 138 -2109 172
rect -2019 138 -1851 172
rect -1761 138 -1593 172
rect -1503 138 -1335 172
rect -1245 138 -1077 172
rect -987 138 -819 172
rect -729 138 -561 172
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect 561 138 729 172
rect 819 138 987 172
rect 1077 138 1245 172
rect 1335 138 1503 172
rect 1593 138 1761 172
rect 1851 138 2019 172
rect 2109 138 2277 172
rect 2367 138 2535 172
rect 2625 138 2793 172
rect 2883 138 3051 172
rect 3141 138 3309 172
rect 3399 138 3567 172
rect 3657 138 3825 172
rect -3825 -172 -3657 -138
rect -3567 -172 -3399 -138
rect -3309 -172 -3141 -138
rect -3051 -172 -2883 -138
rect -2793 -172 -2625 -138
rect -2535 -172 -2367 -138
rect -2277 -172 -2109 -138
rect -2019 -172 -1851 -138
rect -1761 -172 -1593 -138
rect -1503 -172 -1335 -138
rect -1245 -172 -1077 -138
rect -987 -172 -819 -138
rect -729 -172 -561 -138
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
rect 561 -172 729 -138
rect 819 -172 987 -138
rect 1077 -172 1245 -138
rect 1335 -172 1503 -138
rect 1593 -172 1761 -138
rect 1851 -172 2019 -138
rect 2109 -172 2277 -138
rect 2367 -172 2535 -138
rect 2625 -172 2793 -138
rect 2883 -172 3051 -138
rect 3141 -172 3309 -138
rect 3399 -172 3567 -138
rect 3657 -172 3825 -138
<< locali >>
rect -4001 240 -3905 274
rect 3905 240 4001 274
rect -4001 178 -3967 240
rect 3967 178 4001 240
rect -3841 138 -3825 172
rect -3657 138 -3641 172
rect -3583 138 -3567 172
rect -3399 138 -3383 172
rect -3325 138 -3309 172
rect -3141 138 -3125 172
rect -3067 138 -3051 172
rect -2883 138 -2867 172
rect -2809 138 -2793 172
rect -2625 138 -2609 172
rect -2551 138 -2535 172
rect -2367 138 -2351 172
rect -2293 138 -2277 172
rect -2109 138 -2093 172
rect -2035 138 -2019 172
rect -1851 138 -1835 172
rect -1777 138 -1761 172
rect -1593 138 -1577 172
rect -1519 138 -1503 172
rect -1335 138 -1319 172
rect -1261 138 -1245 172
rect -1077 138 -1061 172
rect -1003 138 -987 172
rect -819 138 -803 172
rect -745 138 -729 172
rect -561 138 -545 172
rect -487 138 -471 172
rect -303 138 -287 172
rect -229 138 -213 172
rect -45 138 -29 172
rect 29 138 45 172
rect 213 138 229 172
rect 287 138 303 172
rect 471 138 487 172
rect 545 138 561 172
rect 729 138 745 172
rect 803 138 819 172
rect 987 138 1003 172
rect 1061 138 1077 172
rect 1245 138 1261 172
rect 1319 138 1335 172
rect 1503 138 1519 172
rect 1577 138 1593 172
rect 1761 138 1777 172
rect 1835 138 1851 172
rect 2019 138 2035 172
rect 2093 138 2109 172
rect 2277 138 2293 172
rect 2351 138 2367 172
rect 2535 138 2551 172
rect 2609 138 2625 172
rect 2793 138 2809 172
rect 2867 138 2883 172
rect 3051 138 3067 172
rect 3125 138 3141 172
rect 3309 138 3325 172
rect 3383 138 3399 172
rect 3567 138 3583 172
rect 3641 138 3657 172
rect 3825 138 3841 172
rect -3887 88 -3853 104
rect -3887 -104 -3853 -88
rect -3629 88 -3595 104
rect -3629 -104 -3595 -88
rect -3371 88 -3337 104
rect -3371 -104 -3337 -88
rect -3113 88 -3079 104
rect -3113 -104 -3079 -88
rect -2855 88 -2821 104
rect -2855 -104 -2821 -88
rect -2597 88 -2563 104
rect -2597 -104 -2563 -88
rect -2339 88 -2305 104
rect -2339 -104 -2305 -88
rect -2081 88 -2047 104
rect -2081 -104 -2047 -88
rect -1823 88 -1789 104
rect -1823 -104 -1789 -88
rect -1565 88 -1531 104
rect -1565 -104 -1531 -88
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect 1531 88 1565 104
rect 1531 -104 1565 -88
rect 1789 88 1823 104
rect 1789 -104 1823 -88
rect 2047 88 2081 104
rect 2047 -104 2081 -88
rect 2305 88 2339 104
rect 2305 -104 2339 -88
rect 2563 88 2597 104
rect 2563 -104 2597 -88
rect 2821 88 2855 104
rect 2821 -104 2855 -88
rect 3079 88 3113 104
rect 3079 -104 3113 -88
rect 3337 88 3371 104
rect 3337 -104 3371 -88
rect 3595 88 3629 104
rect 3595 -104 3629 -88
rect 3853 88 3887 104
rect 3853 -104 3887 -88
rect -3841 -172 -3825 -138
rect -3657 -172 -3641 -138
rect -3583 -172 -3567 -138
rect -3399 -172 -3383 -138
rect -3325 -172 -3309 -138
rect -3141 -172 -3125 -138
rect -3067 -172 -3051 -138
rect -2883 -172 -2867 -138
rect -2809 -172 -2793 -138
rect -2625 -172 -2609 -138
rect -2551 -172 -2535 -138
rect -2367 -172 -2351 -138
rect -2293 -172 -2277 -138
rect -2109 -172 -2093 -138
rect -2035 -172 -2019 -138
rect -1851 -172 -1835 -138
rect -1777 -172 -1761 -138
rect -1593 -172 -1577 -138
rect -1519 -172 -1503 -138
rect -1335 -172 -1319 -138
rect -1261 -172 -1245 -138
rect -1077 -172 -1061 -138
rect -1003 -172 -987 -138
rect -819 -172 -803 -138
rect -745 -172 -729 -138
rect -561 -172 -545 -138
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 545 -172 561 -138
rect 729 -172 745 -138
rect 803 -172 819 -138
rect 987 -172 1003 -138
rect 1061 -172 1077 -138
rect 1245 -172 1261 -138
rect 1319 -172 1335 -138
rect 1503 -172 1519 -138
rect 1577 -172 1593 -138
rect 1761 -172 1777 -138
rect 1835 -172 1851 -138
rect 2019 -172 2035 -138
rect 2093 -172 2109 -138
rect 2277 -172 2293 -138
rect 2351 -172 2367 -138
rect 2535 -172 2551 -138
rect 2609 -172 2625 -138
rect 2793 -172 2809 -138
rect 2867 -172 2883 -138
rect 3051 -172 3067 -138
rect 3125 -172 3141 -138
rect 3309 -172 3325 -138
rect 3383 -172 3399 -138
rect 3567 -172 3583 -138
rect 3641 -172 3657 -138
rect 3825 -172 3841 -138
rect -4001 -240 -3967 -178
rect 3967 -240 4001 -178
rect -4001 -274 -3905 -240
rect 3905 -274 4001 -240
<< viali >>
rect -3825 138 -3657 172
rect -3567 138 -3399 172
rect -3309 138 -3141 172
rect -3051 138 -2883 172
rect -2793 138 -2625 172
rect -2535 138 -2367 172
rect -2277 138 -2109 172
rect -2019 138 -1851 172
rect -1761 138 -1593 172
rect -1503 138 -1335 172
rect -1245 138 -1077 172
rect -987 138 -819 172
rect -729 138 -561 172
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect 561 138 729 172
rect 819 138 987 172
rect 1077 138 1245 172
rect 1335 138 1503 172
rect 1593 138 1761 172
rect 1851 138 2019 172
rect 2109 138 2277 172
rect 2367 138 2535 172
rect 2625 138 2793 172
rect 2883 138 3051 172
rect 3141 138 3309 172
rect 3399 138 3567 172
rect 3657 138 3825 172
rect -3887 -88 -3853 88
rect -3629 -88 -3595 88
rect -3371 -88 -3337 88
rect -3113 -88 -3079 88
rect -2855 -88 -2821 88
rect -2597 -88 -2563 88
rect -2339 -88 -2305 88
rect -2081 -88 -2047 88
rect -1823 -88 -1789 88
rect -1565 -88 -1531 88
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect 1531 -88 1565 88
rect 1789 -88 1823 88
rect 2047 -88 2081 88
rect 2305 -88 2339 88
rect 2563 -88 2597 88
rect 2821 -88 2855 88
rect 3079 -88 3113 88
rect 3337 -88 3371 88
rect 3595 -88 3629 88
rect 3853 -88 3887 88
rect -3825 -172 -3657 -138
rect -3567 -172 -3399 -138
rect -3309 -172 -3141 -138
rect -3051 -172 -2883 -138
rect -2793 -172 -2625 -138
rect -2535 -172 -2367 -138
rect -2277 -172 -2109 -138
rect -2019 -172 -1851 -138
rect -1761 -172 -1593 -138
rect -1503 -172 -1335 -138
rect -1245 -172 -1077 -138
rect -987 -172 -819 -138
rect -729 -172 -561 -138
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
rect 561 -172 729 -138
rect 819 -172 987 -138
rect 1077 -172 1245 -138
rect 1335 -172 1503 -138
rect 1593 -172 1761 -138
rect 1851 -172 2019 -138
rect 2109 -172 2277 -138
rect 2367 -172 2535 -138
rect 2625 -172 2793 -138
rect 2883 -172 3051 -138
rect 3141 -172 3309 -138
rect 3399 -172 3567 -138
rect 3657 -172 3825 -138
<< metal1 >>
rect -3837 172 -3645 178
rect -3837 138 -3825 172
rect -3657 138 -3645 172
rect -3837 132 -3645 138
rect -3579 172 -3387 178
rect -3579 138 -3567 172
rect -3399 138 -3387 172
rect -3579 132 -3387 138
rect -3321 172 -3129 178
rect -3321 138 -3309 172
rect -3141 138 -3129 172
rect -3321 132 -3129 138
rect -3063 172 -2871 178
rect -3063 138 -3051 172
rect -2883 138 -2871 172
rect -3063 132 -2871 138
rect -2805 172 -2613 178
rect -2805 138 -2793 172
rect -2625 138 -2613 172
rect -2805 132 -2613 138
rect -2547 172 -2355 178
rect -2547 138 -2535 172
rect -2367 138 -2355 172
rect -2547 132 -2355 138
rect -2289 172 -2097 178
rect -2289 138 -2277 172
rect -2109 138 -2097 172
rect -2289 132 -2097 138
rect -2031 172 -1839 178
rect -2031 138 -2019 172
rect -1851 138 -1839 172
rect -2031 132 -1839 138
rect -1773 172 -1581 178
rect -1773 138 -1761 172
rect -1593 138 -1581 172
rect -1773 132 -1581 138
rect -1515 172 -1323 178
rect -1515 138 -1503 172
rect -1335 138 -1323 172
rect -1515 132 -1323 138
rect -1257 172 -1065 178
rect -1257 138 -1245 172
rect -1077 138 -1065 172
rect -1257 132 -1065 138
rect -999 172 -807 178
rect -999 138 -987 172
rect -819 138 -807 172
rect -999 132 -807 138
rect -741 172 -549 178
rect -741 138 -729 172
rect -561 138 -549 172
rect -741 132 -549 138
rect -483 172 -291 178
rect -483 138 -471 172
rect -303 138 -291 172
rect -483 132 -291 138
rect -225 172 -33 178
rect -225 138 -213 172
rect -45 138 -33 172
rect -225 132 -33 138
rect 33 172 225 178
rect 33 138 45 172
rect 213 138 225 172
rect 33 132 225 138
rect 291 172 483 178
rect 291 138 303 172
rect 471 138 483 172
rect 291 132 483 138
rect 549 172 741 178
rect 549 138 561 172
rect 729 138 741 172
rect 549 132 741 138
rect 807 172 999 178
rect 807 138 819 172
rect 987 138 999 172
rect 807 132 999 138
rect 1065 172 1257 178
rect 1065 138 1077 172
rect 1245 138 1257 172
rect 1065 132 1257 138
rect 1323 172 1515 178
rect 1323 138 1335 172
rect 1503 138 1515 172
rect 1323 132 1515 138
rect 1581 172 1773 178
rect 1581 138 1593 172
rect 1761 138 1773 172
rect 1581 132 1773 138
rect 1839 172 2031 178
rect 1839 138 1851 172
rect 2019 138 2031 172
rect 1839 132 2031 138
rect 2097 172 2289 178
rect 2097 138 2109 172
rect 2277 138 2289 172
rect 2097 132 2289 138
rect 2355 172 2547 178
rect 2355 138 2367 172
rect 2535 138 2547 172
rect 2355 132 2547 138
rect 2613 172 2805 178
rect 2613 138 2625 172
rect 2793 138 2805 172
rect 2613 132 2805 138
rect 2871 172 3063 178
rect 2871 138 2883 172
rect 3051 138 3063 172
rect 2871 132 3063 138
rect 3129 172 3321 178
rect 3129 138 3141 172
rect 3309 138 3321 172
rect 3129 132 3321 138
rect 3387 172 3579 178
rect 3387 138 3399 172
rect 3567 138 3579 172
rect 3387 132 3579 138
rect 3645 172 3837 178
rect 3645 138 3657 172
rect 3825 138 3837 172
rect 3645 132 3837 138
rect -3893 88 -3847 100
rect -3893 -88 -3887 88
rect -3853 -88 -3847 88
rect -3893 -100 -3847 -88
rect -3635 88 -3589 100
rect -3635 -88 -3629 88
rect -3595 -88 -3589 88
rect -3635 -100 -3589 -88
rect -3377 88 -3331 100
rect -3377 -88 -3371 88
rect -3337 -88 -3331 88
rect -3377 -100 -3331 -88
rect -3119 88 -3073 100
rect -3119 -88 -3113 88
rect -3079 -88 -3073 88
rect -3119 -100 -3073 -88
rect -2861 88 -2815 100
rect -2861 -88 -2855 88
rect -2821 -88 -2815 88
rect -2861 -100 -2815 -88
rect -2603 88 -2557 100
rect -2603 -88 -2597 88
rect -2563 -88 -2557 88
rect -2603 -100 -2557 -88
rect -2345 88 -2299 100
rect -2345 -88 -2339 88
rect -2305 -88 -2299 88
rect -2345 -100 -2299 -88
rect -2087 88 -2041 100
rect -2087 -88 -2081 88
rect -2047 -88 -2041 88
rect -2087 -100 -2041 -88
rect -1829 88 -1783 100
rect -1829 -88 -1823 88
rect -1789 -88 -1783 88
rect -1829 -100 -1783 -88
rect -1571 88 -1525 100
rect -1571 -88 -1565 88
rect -1531 -88 -1525 88
rect -1571 -100 -1525 -88
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect 1525 88 1571 100
rect 1525 -88 1531 88
rect 1565 -88 1571 88
rect 1525 -100 1571 -88
rect 1783 88 1829 100
rect 1783 -88 1789 88
rect 1823 -88 1829 88
rect 1783 -100 1829 -88
rect 2041 88 2087 100
rect 2041 -88 2047 88
rect 2081 -88 2087 88
rect 2041 -100 2087 -88
rect 2299 88 2345 100
rect 2299 -88 2305 88
rect 2339 -88 2345 88
rect 2299 -100 2345 -88
rect 2557 88 2603 100
rect 2557 -88 2563 88
rect 2597 -88 2603 88
rect 2557 -100 2603 -88
rect 2815 88 2861 100
rect 2815 -88 2821 88
rect 2855 -88 2861 88
rect 2815 -100 2861 -88
rect 3073 88 3119 100
rect 3073 -88 3079 88
rect 3113 -88 3119 88
rect 3073 -100 3119 -88
rect 3331 88 3377 100
rect 3331 -88 3337 88
rect 3371 -88 3377 88
rect 3331 -100 3377 -88
rect 3589 88 3635 100
rect 3589 -88 3595 88
rect 3629 -88 3635 88
rect 3589 -100 3635 -88
rect 3847 88 3893 100
rect 3847 -88 3853 88
rect 3887 -88 3893 88
rect 3847 -100 3893 -88
rect -3837 -138 -3645 -132
rect -3837 -172 -3825 -138
rect -3657 -172 -3645 -138
rect -3837 -178 -3645 -172
rect -3579 -138 -3387 -132
rect -3579 -172 -3567 -138
rect -3399 -172 -3387 -138
rect -3579 -178 -3387 -172
rect -3321 -138 -3129 -132
rect -3321 -172 -3309 -138
rect -3141 -172 -3129 -138
rect -3321 -178 -3129 -172
rect -3063 -138 -2871 -132
rect -3063 -172 -3051 -138
rect -2883 -172 -2871 -138
rect -3063 -178 -2871 -172
rect -2805 -138 -2613 -132
rect -2805 -172 -2793 -138
rect -2625 -172 -2613 -138
rect -2805 -178 -2613 -172
rect -2547 -138 -2355 -132
rect -2547 -172 -2535 -138
rect -2367 -172 -2355 -138
rect -2547 -178 -2355 -172
rect -2289 -138 -2097 -132
rect -2289 -172 -2277 -138
rect -2109 -172 -2097 -138
rect -2289 -178 -2097 -172
rect -2031 -138 -1839 -132
rect -2031 -172 -2019 -138
rect -1851 -172 -1839 -138
rect -2031 -178 -1839 -172
rect -1773 -138 -1581 -132
rect -1773 -172 -1761 -138
rect -1593 -172 -1581 -138
rect -1773 -178 -1581 -172
rect -1515 -138 -1323 -132
rect -1515 -172 -1503 -138
rect -1335 -172 -1323 -138
rect -1515 -178 -1323 -172
rect -1257 -138 -1065 -132
rect -1257 -172 -1245 -138
rect -1077 -172 -1065 -138
rect -1257 -178 -1065 -172
rect -999 -138 -807 -132
rect -999 -172 -987 -138
rect -819 -172 -807 -138
rect -999 -178 -807 -172
rect -741 -138 -549 -132
rect -741 -172 -729 -138
rect -561 -172 -549 -138
rect -741 -178 -549 -172
rect -483 -138 -291 -132
rect -483 -172 -471 -138
rect -303 -172 -291 -138
rect -483 -178 -291 -172
rect -225 -138 -33 -132
rect -225 -172 -213 -138
rect -45 -172 -33 -138
rect -225 -178 -33 -172
rect 33 -138 225 -132
rect 33 -172 45 -138
rect 213 -172 225 -138
rect 33 -178 225 -172
rect 291 -138 483 -132
rect 291 -172 303 -138
rect 471 -172 483 -138
rect 291 -178 483 -172
rect 549 -138 741 -132
rect 549 -172 561 -138
rect 729 -172 741 -138
rect 549 -178 741 -172
rect 807 -138 999 -132
rect 807 -172 819 -138
rect 987 -172 999 -138
rect 807 -178 999 -172
rect 1065 -138 1257 -132
rect 1065 -172 1077 -138
rect 1245 -172 1257 -138
rect 1065 -178 1257 -172
rect 1323 -138 1515 -132
rect 1323 -172 1335 -138
rect 1503 -172 1515 -138
rect 1323 -178 1515 -172
rect 1581 -138 1773 -132
rect 1581 -172 1593 -138
rect 1761 -172 1773 -138
rect 1581 -178 1773 -172
rect 1839 -138 2031 -132
rect 1839 -172 1851 -138
rect 2019 -172 2031 -138
rect 1839 -178 2031 -172
rect 2097 -138 2289 -132
rect 2097 -172 2109 -138
rect 2277 -172 2289 -138
rect 2097 -178 2289 -172
rect 2355 -138 2547 -132
rect 2355 -172 2367 -138
rect 2535 -172 2547 -138
rect 2355 -178 2547 -172
rect 2613 -138 2805 -132
rect 2613 -172 2625 -138
rect 2793 -172 2805 -138
rect 2613 -178 2805 -172
rect 2871 -138 3063 -132
rect 2871 -172 2883 -138
rect 3051 -172 3063 -138
rect 2871 -178 3063 -172
rect 3129 -138 3321 -132
rect 3129 -172 3141 -138
rect 3309 -172 3321 -138
rect 3129 -178 3321 -172
rect 3387 -138 3579 -132
rect 3387 -172 3399 -138
rect 3567 -172 3579 -138
rect 3387 -178 3579 -172
rect 3645 -138 3837 -132
rect 3645 -172 3657 -138
rect 3825 -172 3837 -138
rect 3645 -178 3837 -172
<< properties >>
string FIXED_BBOX -3984 -257 3984 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
