magic
tech sky130A
magscale 1 2
timestamp 1698088655
<< locali >>
rect -15648 68202 -15148 69252
rect -16698 67702 -15148 68202
rect -15648 67652 -15148 67702
rect -15098 67652 -14598 69252
rect -16698 67152 -14598 67652
rect -15098 67102 -14598 67152
rect -14548 67102 -14048 69252
rect -16698 66602 -14048 67102
rect -14548 66552 -14048 66602
rect -13998 66552 -13498 69252
rect -16698 66052 -13498 66552
rect -13998 66002 -13498 66052
rect -13448 66002 -12948 69252
rect -16698 65502 -12948 66002
rect -13448 65452 -12948 65502
rect -12898 65452 -12398 69252
rect -16698 64952 -12398 65452
rect -12898 64902 -12398 64952
rect -12348 64902 -11848 69252
rect -16698 64402 -11848 64902
rect -12348 64352 -11848 64402
rect -11798 64352 -11298 69252
rect -16698 63852 -11298 64352
rect -11798 63802 -11298 63852
rect -11248 63802 -10748 69252
rect -16698 63302 -10748 63802
rect -11248 63252 -10748 63302
rect -10698 63252 -10198 69252
rect -16698 62752 -10198 63252
rect -10698 62702 -10198 62752
rect -10148 62702 -9648 69252
rect -16698 62202 -9648 62702
rect -10148 62152 -9648 62202
rect -9598 62152 -9098 69252
rect -16698 61652 -9098 62152
rect -9598 61602 -9098 61652
rect -9048 61602 -8548 69252
rect -16698 61102 -8548 61602
rect -9048 61052 -8548 61102
rect -8498 61052 -7998 69252
rect -16698 60552 -7998 61052
rect -8498 60502 -7998 60552
rect -7948 60502 -7448 69252
rect -16698 60002 -7448 60502
rect -7948 59952 -7448 60002
rect -7398 59952 -6898 69252
rect -16698 59452 -6898 59952
rect -7398 59402 -6898 59452
rect -6848 59402 -6348 69252
rect -16698 58902 -6348 59402
rect -6848 58852 -6348 58902
rect -6298 58852 -5798 69252
rect -16698 58352 -5798 58852
rect -6298 58302 -5798 58352
rect -5748 58302 -5248 69252
rect -16698 57802 -5248 58302
rect -5748 57752 -5248 57802
rect -5198 57752 -4698 69252
rect -16698 57252 -4698 57752
rect -5198 57202 -4698 57252
rect -4648 57202 -4148 69252
rect -16698 56702 -4148 57202
rect -4648 56652 -4148 56702
rect -4098 56652 -3598 69252
rect -16698 56152 -3598 56652
rect -4098 56102 -3598 56152
rect -3548 56102 -3048 69252
rect -16698 55602 -3048 56102
rect -3548 55552 -3048 55602
rect -2998 55552 -2498 69252
rect -16698 55052 -2498 55552
rect -2998 55002 -2498 55052
rect -2448 55002 -1948 69252
rect -16698 54502 -1948 55002
rect -2448 54452 -1948 54502
rect -1898 54452 -1398 69252
rect -16698 53952 -1398 54452
rect -1898 53902 -1398 53952
rect -1348 53902 -848 69252
rect -16698 53402 -848 53902
rect -1348 53352 -848 53402
rect -798 53352 -298 69252
rect -16698 52852 -298 53352
rect -798 52802 -298 52852
rect -248 52802 252 69252
rect 302 53352 802 69252
rect 852 53902 1352 69252
rect 1402 54452 1902 69252
rect 1952 55002 2452 69252
rect 2502 55552 3002 69252
rect 3052 56102 3552 69252
rect 3602 56652 4102 69252
rect 4152 57202 4652 69252
rect 4702 57752 5202 69252
rect 5252 58302 5752 69252
rect 5802 58852 6302 69252
rect 6352 59402 6852 69252
rect 6902 59952 7402 69252
rect 7452 60502 7952 69252
rect 8002 61052 8502 69252
rect 8552 61602 9052 69252
rect 9102 62152 9602 69252
rect 9652 62702 10152 69252
rect 10202 63252 10702 69252
rect 10752 63802 11252 69252
rect 11302 64352 11802 69252
rect 11852 64902 12352 69252
rect 12402 65452 12902 69252
rect 12952 66002 13452 69252
rect 13502 66552 14002 69252
rect 14052 67102 14552 69252
rect 14602 67652 15102 69252
rect 15152 68202 15652 69252
rect 15152 67702 16702 68202
rect 15152 67652 15652 67702
rect 14602 67152 16702 67652
rect 14602 67102 15102 67152
rect 14052 66602 16702 67102
rect 14052 66552 14552 66602
rect 13502 66052 16702 66552
rect 13502 66002 14002 66052
rect 12952 65502 16702 66002
rect 12952 65452 13452 65502
rect 12402 64952 16702 65452
rect 12402 64902 12902 64952
rect 11852 64402 16702 64902
rect 11852 64352 12352 64402
rect 11302 63852 16702 64352
rect 11302 63802 11802 63852
rect 10752 63302 16702 63802
rect 10752 63252 11252 63302
rect 10202 62752 16702 63252
rect 10202 62702 10702 62752
rect 9652 62202 16702 62702
rect 9652 62152 10152 62202
rect 9102 61652 16702 62152
rect 9102 61602 9602 61652
rect 8552 61102 16702 61602
rect 8552 61052 9052 61102
rect 8002 60552 16702 61052
rect 8002 60502 8502 60552
rect 7452 60002 16702 60502
rect 7452 59952 7952 60002
rect 6902 59452 16702 59952
rect 6902 59402 7402 59452
rect 6352 58902 16702 59402
rect 6352 58852 6852 58902
rect 5802 58352 16702 58852
rect 5802 58302 6302 58352
rect 5252 57802 16702 58302
rect 5252 57752 5752 57802
rect 4702 57252 16702 57752
rect 4702 57202 5202 57252
rect 4152 56702 16702 57202
rect 4152 56652 4652 56702
rect 3602 56152 16702 56652
rect 3602 56102 4102 56152
rect 3052 55602 16702 56102
rect 3052 55552 3552 55602
rect 2502 55052 16702 55552
rect 2502 55002 3002 55052
rect 1952 54502 16702 55002
rect 1952 54452 2452 54502
rect 1402 53952 16702 54452
rect 1402 53902 1902 53952
rect 852 53402 16702 53902
rect 852 53352 1352 53402
rect 302 52852 16702 53352
rect 302 52802 802 52852
rect -16698 52783 16702 52802
rect -16698 52302 -224 52783
rect -248 52252 -224 52302
rect -16698 51752 -224 52252
rect -248 51702 -224 51752
rect -16698 51223 -224 51702
rect 236 52302 16702 52783
rect 236 52252 252 52302
rect 236 51752 16702 52252
rect 236 51702 252 51752
rect 236 51223 16702 51702
rect -16698 51202 16702 51223
rect -798 51152 -298 51202
rect -16698 50652 -298 51152
rect -1348 50602 -848 50652
rect -16698 50102 -848 50602
rect -1898 50052 -1398 50102
rect -16698 49552 -1398 50052
rect -2448 49502 -1948 49552
rect -16698 49002 -1948 49502
rect -2998 48952 -2498 49002
rect -16698 48452 -2498 48952
rect -3548 48402 -3048 48452
rect -16698 47902 -3048 48402
rect -4098 47852 -3598 47902
rect -16698 47352 -3598 47852
rect -4648 47302 -4148 47352
rect -16698 46802 -4148 47302
rect -5198 46752 -4698 46802
rect -16698 46252 -4698 46752
rect -5748 46202 -5248 46252
rect -16698 45702 -5248 46202
rect -6298 45652 -5798 45702
rect -16698 45152 -5798 45652
rect -6848 45102 -6348 45152
rect -16698 44602 -6348 45102
rect -7398 44552 -6898 44602
rect -16698 44052 -6898 44552
rect -7948 44002 -7448 44052
rect -16698 43502 -7448 44002
rect -8498 43452 -7998 43502
rect -16698 42952 -7998 43452
rect -9048 42902 -8548 42952
rect -16698 42402 -8548 42902
rect -9598 42352 -9098 42402
rect -16698 41852 -9098 42352
rect -10148 41802 -9648 41852
rect -16698 41302 -9648 41802
rect -10698 41252 -10198 41302
rect -16698 40752 -10198 41252
rect -11248 40702 -10748 40752
rect -16698 40202 -10748 40702
rect -11798 40152 -11298 40202
rect -16698 39652 -11298 40152
rect -12348 39602 -11848 39652
rect -16698 39102 -11848 39602
rect -12898 39052 -12398 39102
rect -16698 38552 -12398 39052
rect -13448 38502 -12948 38552
rect -16698 38002 -12948 38502
rect -13998 37952 -13498 38002
rect -16698 37452 -13498 37952
rect -14548 37402 -14048 37452
rect -16698 36902 -14048 37402
rect -15098 36852 -14598 36902
rect -16698 36352 -14598 36852
rect -15648 35352 -15148 36352
rect -15098 35352 -14598 36352
rect -14548 35352 -14048 36902
rect -13998 35352 -13498 37452
rect -13448 35352 -12948 38002
rect -12898 35352 -12398 38552
rect -12348 35352 -11848 39102
rect -11798 35352 -11298 39652
rect -11248 35352 -10748 40202
rect -10698 35352 -10198 40752
rect -10148 35352 -9648 41302
rect -9598 35352 -9098 41852
rect -9048 35352 -8548 42402
rect -8498 35352 -7998 42952
rect -7948 35352 -7448 43502
rect -7398 35352 -6898 44052
rect -6848 35352 -6348 44602
rect -6298 35352 -5798 45152
rect -5748 35352 -5248 45702
rect -5198 35352 -4698 46252
rect -4648 35352 -4148 46802
rect -4098 35352 -3598 47352
rect -3548 35352 -3048 47902
rect -2998 35352 -2498 48452
rect -2448 35352 -1948 49002
rect -1898 35352 -1398 49552
rect -1348 35352 -848 50102
rect -798 35352 -298 50652
rect -248 35352 252 51202
rect 302 51152 802 51202
rect 302 50652 16702 51152
rect 302 35352 802 50652
rect 852 50602 1352 50652
rect 852 50102 16702 50602
rect 852 35352 1352 50102
rect 1402 50052 1902 50102
rect 1402 49552 16702 50052
rect 1402 35352 1902 49552
rect 1952 49502 2452 49552
rect 1952 49002 16702 49502
rect 1952 35352 2452 49002
rect 2502 48952 3002 49002
rect 2502 48452 16702 48952
rect 2502 35352 3002 48452
rect 3052 48402 3552 48452
rect 3052 47902 16702 48402
rect 3052 35352 3552 47902
rect 3602 47852 4102 47902
rect 3602 47352 16702 47852
rect 3602 35352 4102 47352
rect 4152 47302 4652 47352
rect 4152 46802 16702 47302
rect 4152 35352 4652 46802
rect 4702 46752 5202 46802
rect 4702 46252 16702 46752
rect 4702 35352 5202 46252
rect 5252 46202 5752 46252
rect 5252 45702 16702 46202
rect 5252 35352 5752 45702
rect 5802 45652 6302 45702
rect 5802 45152 16702 45652
rect 5802 35352 6302 45152
rect 6352 45102 6852 45152
rect 6352 44602 16702 45102
rect 6352 35352 6852 44602
rect 6902 44552 7402 44602
rect 6902 44052 16702 44552
rect 6902 35352 7402 44052
rect 7452 44002 7952 44052
rect 7452 43502 16702 44002
rect 7452 35352 7952 43502
rect 8002 43452 8502 43502
rect 8002 42952 16702 43452
rect 8002 35352 8502 42952
rect 8552 42902 9052 42952
rect 8552 42402 16702 42902
rect 8552 35352 9052 42402
rect 9102 42352 9602 42402
rect 9102 41852 16702 42352
rect 9102 35352 9602 41852
rect 9652 41802 10152 41852
rect 9652 41302 16702 41802
rect 9652 35352 10152 41302
rect 10202 41252 10702 41302
rect 10202 40752 16702 41252
rect 10202 35352 10702 40752
rect 10752 40702 11252 40752
rect 10752 40202 16702 40702
rect 10752 35352 11252 40202
rect 11302 40152 11802 40202
rect 11302 39652 16702 40152
rect 11302 35352 11802 39652
rect 11852 39602 12352 39652
rect 11852 39102 16702 39602
rect 11852 35352 12352 39102
rect 12402 39052 12902 39102
rect 12402 38552 16702 39052
rect 12402 35352 12902 38552
rect 12952 38502 13452 38552
rect 12952 38002 16702 38502
rect 12952 35352 13452 38002
rect 13502 37952 14002 38002
rect 13502 37452 16702 37952
rect 13502 35352 14002 37452
rect 14052 37402 14552 37452
rect 14052 36902 16702 37402
rect 14052 35352 14552 36902
rect 14602 36852 15102 36902
rect 14602 36352 16702 36852
rect 14602 35352 15102 36352
rect 15152 35352 15652 36352
<< viali >>
rect -224 51223 236 52783
<< metal1 >>
rect -244 52783 16756 52803
rect -244 51223 -224 52783
rect 236 51223 16756 52783
rect -244 51203 16756 51223
<< metal4 >>
rect -6620 68400 -1793 68500
rect -6620 67600 -6527 68400
rect -2600 67784 -1793 68400
tri -1793 67784 -1077 68500 sw
rect -2600 67600 -1077 67784
rect -6620 67500 -1077 67600
tri -2207 66500 -1207 67500 ne
rect -1207 66586 -1077 67500
tri -1077 66586 121 67784 sw
rect -1207 66500 121 66586
rect -5210 66400 -2163 66500
rect -5210 65600 -5110 66400
rect -2600 65630 -2163 66400
tri -2163 65630 -1293 66500 sw
tri -1207 65630 -337 66500 ne
rect -337 65630 121 66500
rect -2600 65600 -1293 65630
rect -5210 65500 -1293 65600
tri -2577 65293 -2370 65500 ne
rect -2370 65414 -1293 65500
tri -1293 65414 -1077 65630 sw
rect -2370 65293 -1077 65414
tri -2370 64000 -1077 65293 ne
tri -1077 65172 -835 65414 sw
tri -337 65172 121 65630 ne
tri 121 65172 1535 66586 sw
rect -1077 64400 -835 65172
tri -835 64400 -63 65172 sw
tri 121 64400 893 65172 ne
rect 893 64500 1535 65172
tri 1535 64500 2207 65172 sw
rect 893 64400 4960 64500
rect -1077 64360 710 64400
rect -1077 64000 -390 64360
tri -1077 63600 -677 64000 ne
rect -677 63640 -390 64000
rect 670 63640 710 64360
rect -677 63600 710 63640
tri 893 63500 1793 64400 ne
rect 1793 63600 2600 64400
rect 4871 63600 4960 64400
rect 1793 63500 4960 63600
rect 15500 58740 16500 58835
rect 11500 57080 12500 57178
rect -10450 56042 -9450 56142
rect -10450 54600 -10350 56042
rect -9550 54600 -9450 56042
tri -11122 53535 -10450 54207 se
rect -10450 53793 -9450 54600
rect -10450 53535 -10250 53793
tri -12536 52121 -11122 53535 se
rect -11122 52993 -10250 53535
tri -10250 52993 -9450 53793 nw
rect 11500 53720 11590 57080
rect 12410 53720 12500 57080
tri -11122 52121 -10250 52993 nw
rect -10250 52570 -9450 52620
tri -13950 50707 -12536 52121 se
rect -12536 51807 -11436 52121
tri -11436 51807 -11122 52121 nw
tri -12536 50707 -11436 51807 nw
tri -14450 50207 -13950 50707 se
rect -13950 50207 -13450 50707
rect -14450 49400 -13450 50207
tri -13450 49793 -12536 50707 nw
tri -11364 50693 -10250 51807 se
rect -10250 51580 -10200 52570
rect -9500 51580 -9450 52570
rect -10250 51193 -9450 51580
rect -10250 50693 -9950 51193
tri -9950 50693 -9450 51193 nw
rect -14450 46301 -14350 49400
rect -13550 46301 -13450 49400
tri -12500 49557 -11364 50693 se
rect -11364 49557 -11243 50693
rect -12500 49400 -11243 49557
tri -11243 49400 -9950 50693 nw
rect 11500 50280 12500 53720
rect -12500 46920 -12410 49400
rect -11590 46920 -11500 49400
tri -11500 49143 -11243 49400 nw
rect -12500 46821 -11500 46920
rect 11500 46920 11590 50280
rect 12410 46920 12500 50280
rect 11500 46821 12500 46920
rect 15500 56500 15590 58740
rect 16410 56500 16500 58740
rect 15500 47500 16500 56500
rect -14450 46201 -13450 46301
rect 15500 45270 15600 47500
rect 16400 45270 16500 47500
rect 15500 45166 16500 45270
<< via4 >>
rect -6527 67600 -2600 68400
rect -5110 65600 -2600 66400
rect -390 63640 670 64360
rect 2600 63600 4871 64400
rect -10350 54600 -9550 56042
rect 11590 53720 12410 57080
rect -10200 51580 -9500 52570
rect -14350 46301 -13550 49400
rect -12410 46920 -11590 49400
rect 11590 46920 12410 50280
rect 15590 56500 16410 58740
rect 15600 45270 16400 47500
<< metal5 >>
tri -8041 67293 -6834 68500 se
rect -6834 68400 -2500 68500
rect -6834 67600 -6527 68400
rect -2600 67600 -2500 68400
rect -6834 67500 -2500 67600
rect -6834 67293 -6627 67500
tri -6627 67293 -6420 67500 nw
tri 586 67293 1793 68500 se
rect 1793 68000 6835 68500
tri 6835 68000 7335 68500 sw
rect 1793 67500 7335 68000
rect 1793 67293 1822 67500
tri -9455 65879 -8041 67293 se
tri -8041 65879 -6627 67293 nw
tri -10869 64465 -9455 65879 se
tri -9455 64465 -8041 65879 nw
tri -6627 65829 -5956 66500 se
rect -5956 66400 -2500 66500
rect -5956 65829 -5110 66400
tri -6880 65576 -6627 65829 se
rect -6627 65600 -5110 65829
rect -2600 65600 -2500 66400
tri -828 65879 586 67293 se
rect 586 67115 1822 67293
tri 1822 67115 2207 67500 nw
tri 586 65879 1822 67115 nw
tri 6420 66585 7335 67500 ne
tri 7335 66585 8750 68000 sw
tri 1822 65879 2443 66500 se
rect 2443 66041 6056 66500
tri 6056 66041 6515 66500 sw
tri 7335 66041 7879 66585 ne
rect 7879 66041 8750 66585
rect 2443 65879 6515 66041
rect -6627 65576 -2500 65600
tri -12283 63051 -10869 64465 se
tri -10869 63051 -9455 64465 nw
tri -8041 64415 -6880 65576 se
rect -6880 65500 -2500 65576
tri -8294 64162 -8041 64415 se
rect -8041 64162 -6880 64415
tri -6880 64162 -5542 65500 nw
tri -2207 64500 -828 65879 se
rect -828 65293 0 65879
tri 0 65293 586 65879 nw
tri 1236 65293 1822 65879 se
rect 1822 65500 6515 65879
rect 1822 65293 1857 65500
rect -828 64500 -793 65293
tri -793 64500 0 65293 nw
tri -13697 61637 -12283 63051 se
tri -12283 61637 -10869 63051 nw
tri -9455 63001 -8294 64162 se
rect -8294 63293 -7749 64162
tri -7749 63293 -6880 64162 nw
tri -5542 64135 -5177 64500 se
rect -5177 64135 -1793 64500
tri -6384 63293 -5542 64135 se
rect -5542 63500 -1793 64135
tri -1793 63500 -793 64500 nw
tri 343 64400 1236 65293 se
rect 1236 64500 1857 65293
tri 1857 64500 2857 65500 nw
tri 5642 64627 6515 65500 ne
tri 6515 65170 7386 66041 sw
tri 7879 65170 8750 66041 ne
tri 8750 65170 10165 66585 sw
rect 6515 64627 7386 65170
tri 7386 64627 7929 65170 sw
tri 8750 64627 9293 65170 ne
rect 9293 64627 10165 65170
rect 1236 64400 1357 64500
rect -430 64360 1357 64400
rect -430 63640 -390 64360
rect 670 64000 1357 64360
tri 1357 64000 1857 64500 nw
rect 2500 64400 5178 64500
rect 670 63640 957 64000
rect -430 63600 957 63640
tri 957 63600 1357 64000 nw
rect 2500 63600 2600 64400
rect 4871 64000 5178 64400
tri 5178 64000 5678 64500 sw
tri 6515 64000 7142 64627 ne
rect 7142 64000 7929 64627
rect 4871 63600 5678 64000
rect 2500 63500 5678 63600
rect -5542 63293 -4970 63500
tri -4970 63293 -4763 63500 nw
tri -9708 62748 -9455 63001 se
rect -9455 62748 -8294 63001
tri -8294 62748 -7749 63293 nw
tri -15111 60223 -13697 61637 se
tri -13697 60223 -12283 61637 nw
tri -10869 61587 -9708 62748 se
rect -9708 61879 -9163 62748
tri -9163 61879 -8294 62748 nw
tri -7749 61928 -6384 63293 se
tri -7798 61879 -7749 61928 se
rect -7749 61879 -6384 61928
tri -6384 61879 -4970 63293 nw
tri 4763 62585 5678 63500 ne
tri 5678 62585 7093 64000 sw
tri 7142 63213 7929 64000 ne
tri 7929 63755 8801 64627 sw
tri 9293 63755 10165 64627 ne
tri 10165 63755 11580 65170 sw
rect 7929 63213 8801 63755
tri 8801 63213 9343 63755 sw
tri 10165 63213 10707 63755 ne
rect 10707 63213 11580 63755
tri 7929 62585 8557 63213 ne
rect 8557 62585 9343 63213
tri -11122 61334 -10869 61587 se
rect -10869 61334 -9708 61587
tri -9708 61334 -9163 61879 nw
tri -16496 58838 -15111 60223 se
rect -16500 58809 -15111 58838
tri -15111 58809 -13697 60223 nw
tri -12283 60173 -11122 61334 se
rect -11122 60465 -10577 61334
tri -10577 60465 -9708 61334 nw
tri -9163 60514 -7798 61879 se
tri -9212 60465 -9163 60514 se
rect -9163 60465 -7798 60514
tri -7798 60465 -6384 61879 nw
tri -4970 61829 -4299 62500 se
rect -4299 61829 4399 62500
tri -5708 61091 -4970 61829 se
rect -4970 61798 4399 61829
tri 4399 61798 5101 62500 sw
tri 5678 61798 6465 62585 ne
rect 6465 61798 7093 62585
rect -4970 61500 5101 61798
rect -4970 61091 -4294 61500
tri -4294 61091 -3885 61500 nw
tri -12536 59920 -12283 60173 se
rect -12283 59920 -11122 60173
tri -11122 59920 -10577 60465 nw
rect -16500 45162 -15500 58809
tri -15500 58420 -15111 58809 nw
tri -13697 58759 -12536 59920 se
rect -12536 58759 -12480 59920
tri -14450 58006 -13697 58759 se
rect -13697 58562 -12480 58759
tri -12480 58562 -11122 59920 nw
tri -10577 59100 -9212 60465 se
tri -11115 58562 -10577 59100 se
rect -10577 59051 -9212 59100
tri -9212 59051 -7798 60465 nw
tri -6384 60415 -5708 61091 se
tri -7122 59677 -6384 60415 se
rect -6384 59677 -5708 60415
tri -5708 59677 -4294 61091 nw
tri 3985 60384 5101 61500 ne
tri 5101 61170 5729 61798 sw
tri 6465 61170 7093 61798 ne
tri 7093 61170 8508 62585 sw
tri 8557 61799 9343 62585 ne
tri 9343 62006 10550 63213 sw
tri 10707 62340 11580 63213 ne
tri 11580 62340 12995 63755 sw
tri 11580 62006 11914 62340 ne
rect 11914 62006 12995 62340
rect 9343 61799 10550 62006
tri 9343 61170 9972 61799 ne
rect 9972 61170 10550 61799
rect 5101 60384 5729 61170
tri 5729 60384 6515 61170 sw
tri 7093 60384 7879 61170 ne
rect 7879 60384 8508 61170
rect -10577 58562 -9701 59051
tri -9701 58562 -9212 59051 nw
tri -7798 59001 -7122 59677 se
rect -13697 58006 -13450 58562
rect -14450 54000 -13450 58006
tri -13450 57592 -12480 58562 nw
tri -11991 57686 -11115 58562 se
rect -11115 57686 -10626 58562
tri -12240 57437 -11991 57686 se
rect -11991 57637 -10626 57686
tri -10626 57637 -9701 58562 nw
tri -8536 58263 -7798 59001 se
rect -7798 58263 -7122 59001
tri -7122 58263 -5708 59677 nw
tri 5101 58970 6515 60384 ne
tri 6515 59755 7144 60384 sw
tri 7879 59755 8508 60384 ne
tri 8508 59755 9923 61170 sw
tri 9972 60592 10550 61170 ne
tri 10550 60925 11631 62006 sw
tri 11914 60925 12995 62006 ne
tri 12995 60925 14410 62340 sw
rect 10550 60627 11631 60925
tri 11631 60627 11929 60925 sw
tri 12995 60627 13293 60925 ne
rect 13293 60627 14410 60925
rect 10550 60592 11929 60627
tri 10550 59755 11387 60592 ne
rect 11387 59755 11929 60592
rect 6515 58970 7144 59755
tri 7144 58970 7929 59755 sw
tri 8508 58970 9293 59755 ne
rect 9293 58970 9923 59755
rect -11991 57437 -11500 57637
tri -12480 57198 -12241 57437 se
rect -12241 57198 -11500 57437
tri -12499 57178 -12480 57197 se
rect -12480 57178 -11500 57198
rect -12500 54443 -11500 57178
tri -11500 56763 -10626 57637 nw
tri -9212 57587 -8536 58263 se
tri -9950 56849 -9212 57587 se
rect -9212 56849 -8536 57587
tri -8536 56849 -7122 58263 nw
tri 6515 57556 7929 58970 ne
tri 7929 58340 8559 58970 sw
tri 9293 58340 9923 58970 ne
tri 9923 58340 11338 59755 sw
tri 11387 59213 11929 59755 ne
tri 11929 59510 13046 60627 sw
tri 13293 59510 14410 60627 ne
tri 14410 59510 15825 60925 sw
rect 11929 59213 13046 59510
tri 11929 58340 12802 59213 ne
rect 12802 58420 13046 59213
tri 13046 58420 14136 59510 sw
tri 14410 58420 15500 59510 ne
rect 15500 58835 15825 59510
tri 15825 58835 16500 59510 sw
rect 15500 58740 16500 58835
rect 12802 58340 14136 58420
rect 7929 57556 8559 58340
tri 8559 57556 9343 58340 sw
tri 9923 57556 10707 58340 ne
rect 10707 57556 11338 58340
tri -10450 56349 -9950 56849 se
rect -9950 56349 -9450 56849
rect -10450 56042 -9450 56349
tri -13450 54000 -13243 54207 sw
rect -14450 53793 -13243 54000
tri -14450 52586 -13243 53793 ne
tri -13243 53720 -12963 54000 sw
tri -12500 53720 -11777 54443 ne
rect -11777 53807 -11500 54443
tri -11500 53807 -10450 54857 sw
rect -10450 54600 -10350 56042
rect -9550 54600 -9450 56042
tri -9450 55935 -8536 56849 nw
tri 7929 56142 9343 57556 ne
tri 9343 56349 10550 57556 sw
tri 10707 56925 11338 57556 ne
tri 11338 57179 12499 58340 sw
tri 12802 57592 13550 58340 ne
rect 13550 58006 14136 58340
tri 14136 58006 14550 58420 sw
rect 11338 57080 12500 57179
rect 11338 56925 11590 57080
tri 11338 56763 11500 56925 ne
rect 9343 56142 10550 56349
tri 9343 55935 9550 56142 ne
rect -10450 54500 -9450 54600
rect -11777 53720 -10450 53807
rect -13243 52586 -12963 53720
tri -12963 52586 -11829 53720 sw
tri -11777 52586 -10643 53720 ne
rect -10643 52807 -10450 53720
tri -10450 52807 -9450 53807 sw
rect -10643 52586 -9450 52807
tri -13243 51172 -11829 52586 ne
tri -11829 51414 -10657 52586 sw
tri -10643 52193 -10250 52586 ne
rect -10250 52570 -9450 52586
rect -10250 51580 -10200 52570
rect -9500 51580 -9450 52570
rect -10250 51530 -9450 51580
rect 9550 52500 10550 56142
rect 11500 53720 11590 56925
rect 12410 53720 12500 57080
rect 13550 55728 14550 58006
rect 15500 56500 15590 58740
rect 16410 56500 16500 58740
rect 15500 56400 16500 56500
rect 13550 54728 16752 55728
rect 17266 54728 17366 55728
rect 11500 53623 12500 53720
rect 9550 51500 16852 52500
rect -11829 51172 -10657 51414
tri -11829 50280 -10937 51172 ne
rect -10937 50280 -10657 51172
tri -10657 50280 -9523 51414 sw
tri -10937 49793 -10450 50280 ne
rect -10450 50207 -9523 50280
tri -9523 50207 -9450 50280 sw
rect -14450 49400 -13450 49500
rect -14450 46301 -14350 49400
rect -13550 46301 -13450 49400
rect -12500 49400 -11500 49500
rect -12500 46920 -12410 49400
rect -11590 46920 -11500 49400
rect -10450 47651 -9450 50207
rect -12500 46863 -11500 46920
tri -11500 46863 -11126 47237 sw
tri -10450 46863 -9662 47651 ne
rect -9662 46920 -9450 47651
tri -9450 46920 -8305 48065 sw
tri 8636 47151 9550 48065 se
rect 9550 47651 10550 51500
rect 9550 47151 9819 47651
rect -9662 46863 -8305 46920
rect -12500 46821 -11126 46863
rect -14450 46201 -13450 46301
tri -13450 46201 -13243 46408 sw
rect -14450 45994 -13243 46201
tri -16497 44490 -15825 45162 ne
rect -15825 44530 -15500 45162
tri -15500 44530 -14450 45580 sw
tri -14450 44787 -13243 45994 ne
tri -13243 45457 -12499 46201 sw
tri -12499 45457 -11135 46821 ne
rect -11135 45457 -11126 46821
tri -11126 45457 -9720 46863 sw
tri -9662 45709 -8508 46863 ne
rect -8508 46444 -8305 46863
tri -8305 46444 -7829 46920 sw
rect -8508 45709 -7829 46444
rect -13243 44787 -12499 45457
tri -12499 44787 -11829 45457 sw
rect -15825 44490 -14450 44530
tri -14450 44490 -14410 44530 sw
tri -13243 44490 -12946 44787 ne
rect -12946 44490 -11829 44787
tri -15825 43075 -14410 44490 ne
tri -14410 43075 -12995 44490 sw
tri -12946 43373 -11829 44490 ne
tri -11829 44216 -11258 44787 sw
tri -11135 44216 -9894 45457 ne
rect -9894 44245 -9720 45457
tri -9720 44245 -8508 45457 sw
tri -8508 45270 -8069 45709 ne
rect -8069 45270 -7829 45709
tri -7829 45270 -6655 46444 sw
tri 7222 45737 8636 47151 se
rect 8636 46920 9819 47151
tri 9819 46920 10550 47651 nw
rect 11500 50280 12500 50377
tri 8636 45737 9819 46920 nw
tri 10626 46363 11500 47237 se
rect 11500 46920 11590 50280
rect 12410 46920 12500 50280
rect 11500 46821 12500 46920
rect 13550 48272 16752 49272
rect 17266 48272 17366 49272
rect 11500 46564 12242 46821
tri 12242 46564 12499 46821 nw
rect 11500 46363 12040 46564
tri 12040 46363 12241 46564 nw
tri 10000 45737 10626 46363 se
tri 6942 45457 7222 45737 se
rect 7222 45457 7848 45737
tri -8069 44245 -7044 45270 ne
rect -7044 44245 -6655 45270
tri -6655 44245 -5630 45270 sw
rect -9894 44216 -8508 44245
rect -11829 43373 -11258 44216
tri -11258 43373 -10415 44216 sw
tri -9894 43373 -9051 44216 ne
rect -9051 43373 -8508 44216
tri -11829 43075 -11531 43373 ne
rect -11531 43075 -10415 43373
tri -14410 41660 -12995 43075 ne
tri -12995 41660 -11580 43075 sw
tri -11531 41959 -10415 43075 ne
tri -10415 42830 -9872 43373 sw
tri -9051 42830 -8508 43373 ne
tri -8508 42830 -7093 44245 sw
tri -7044 42879 -5678 44245 ne
rect -5678 43616 -5630 44245
tri -5630 43616 -5001 44245 sw
tri 5701 44216 6942 45457 se
rect 6942 44949 7848 45457
tri 7848 44949 8636 45737 nw
tri 9212 44949 10000 45737 se
rect 10000 44949 10626 45737
tri 10626 44949 12040 46363 nw
tri 12636 45494 13550 46408 se
rect 13550 45994 14550 48272
rect 13550 45494 13747 45994
rect 6942 44323 7222 44949
tri 7222 44323 7848 44949 nw
rect 6942 44216 7115 44323
tri 7115 44216 7222 44323 nw
tri 8479 44216 9212 44949 se
rect -5678 42879 -5001 43616
rect -10415 41959 -9872 42830
tri -9872 41959 -9001 42830 sw
tri -8508 41959 -7637 42830 ne
rect -7637 41959 -7093 42830
tri -10415 41660 -10116 41959 ne
rect -10116 41660 -9001 41959
tri -12995 40245 -11580 41660 ne
tri -11580 40245 -10165 41660 sw
tri -10116 40545 -9001 41660 ne
tri -9001 41415 -8457 41959 sw
tri -7637 41415 -7093 41959 ne
tri -7093 41415 -5678 42830 sw
tri -5678 42202 -5001 42879 ne
tri -5001 42500 -3885 43616 sw
tri 4394 42909 5701 44216 se
rect 5701 42909 5808 44216
tri 5808 42909 7115 44216 nw
tri 7798 43535 8479 44216 se
rect 8479 43535 9212 44216
tri 9212 43535 10626 44949 nw
tri 12040 44898 12636 45494 se
rect 12636 45191 13747 45494
tri 13747 45191 14550 45994 nw
rect 15500 47500 16500 47600
tri 15111 45191 15500 45580 se
rect 15500 45270 15600 47500
rect 16400 45270 16500 47500
rect 15500 45191 16500 45270
tri 11222 44080 12040 44898 se
rect 12040 44080 12636 44898
tri 12636 44080 13747 45191 nw
tri 7172 42909 7798 43535 se
tri 3985 42500 4394 42909 se
rect 4394 42500 5020 42909
rect -5001 42202 5020 42500
tri -5001 41500 -4299 42202 ne
rect -4299 42121 5020 42202
tri 5020 42121 5808 42909 nw
tri 6384 42121 7172 42909 se
rect 7172 42121 7798 42909
tri 7798 42121 9212 43535 nw
tri 10626 43484 11222 44080 se
rect 11222 43777 12333 44080
tri 12333 43777 12636 44080 nw
tri 13747 43827 15111 45191 se
rect 15111 45166 16500 45191
tri 13697 43777 13747 43827 se
rect 13747 43777 15111 43827
tri 15111 43777 16500 45166 nw
tri 9808 42666 10626 43484 se
rect 10626 42666 11222 43484
tri 11222 42666 12333 43777 nw
rect -4299 41500 4399 42121
tri 4399 41500 5020 42121 nw
rect -9001 40545 -8457 41415
tri -8457 40545 -7587 41415 sw
tri -7093 40545 -6223 41415 ne
rect -6223 40545 -5678 41415
tri -9001 40245 -8701 40545 ne
rect -8701 40245 -7587 40545
tri -11580 38830 -10165 40245 ne
tri -10165 38830 -8750 40245 sw
tri -8701 39131 -7587 40245 ne
tri -7587 39242 -6284 40545 sw
tri -6223 40000 -5678 40545 ne
tri -5678 40500 -4763 41415 sw
tri 5020 40757 6384 42121 se
tri 4763 40500 5020 40757 se
rect 5020 40707 6384 40757
tri 6384 40707 7798 42121 nw
tri 9212 42070 9808 42666 se
rect 9808 42363 10919 42666
tri 10919 42363 11222 42666 nw
tri 12333 42413 13697 43777 se
tri 12283 42363 12333 42413 se
rect 12333 42363 13697 42413
tri 13697 42363 15111 43777 nw
tri 8394 41252 9212 42070 se
rect 9212 41252 9808 42070
tri 9808 41252 10919 42363 nw
rect 5020 40500 5177 40707
rect -5678 40000 5177 40500
tri -5678 39500 -5178 40000 ne
rect -5178 39500 5177 40000
tri 5177 39500 6384 40707 nw
tri 7798 40656 8394 41252 se
rect 8394 40949 9505 41252
tri 9505 40949 9808 41252 nw
tri 10919 40999 12283 42363 se
tri 10869 40949 10919 40999 se
rect 10919 40949 12283 40999
tri 12283 40949 13697 42363 nw
tri 6980 39838 7798 40656 se
rect 7798 39838 8394 40656
tri 8394 39838 9505 40949 nw
tri 6384 39242 6980 39838 se
rect 6980 39535 8091 39838
tri 8091 39535 8394 39838 nw
tri 9505 39585 10869 40949 se
tri 9455 39535 9505 39585 se
rect 9505 39535 10869 39585
tri 10869 39535 12283 40949 nw
rect -7587 39131 -6284 39242
tri -6284 39131 -6173 39242 sw
tri -7587 38830 -7286 39131 ne
rect -7286 38830 -6173 39131
tri -10165 37415 -8750 38830 ne
tri -8750 37415 -7335 38830 sw
tri -7286 37717 -6173 38830 ne
tri -6173 38500 -5542 39131 sw
tri 5642 38500 6384 39242 se
rect 6384 38500 6980 39242
rect -6173 38424 6980 38500
tri 6980 38424 8091 39535 nw
rect -6173 37717 6056 38424
tri -6173 37500 -5956 37717 ne
rect -5956 37500 6056 37717
tri 6056 37500 6980 38424 nw
tri 8091 38171 9455 39535 se
tri 8041 38121 8091 38171 se
rect 8091 38121 9455 38171
tri 9455 38121 10869 39535 nw
tri -8750 36000 -7335 37415 ne
tri -7335 36500 -6420 37415 sw
tri 6980 37060 8041 38121 se
tri 6627 36707 6980 37060 se
rect 6980 36707 8041 37060
tri 8041 36707 9455 38121 nw
tri 6420 36500 6627 36707 se
rect 6627 36500 6834 36707
rect -7335 36000 -5427 36500
tri -7335 35500 -6835 36000 ne
rect -6835 35500 -5427 36000
rect -6427 34500 -5427 35500
rect 5427 35500 6834 36500
tri 6834 35500 8041 36707 nw
rect 5427 34500 6427 35500
rect -6427 33886 -5427 33986
rect 5427 33886 6427 33986
use sky130_fd_pr__res_generic_m5_EGUVWD  sky130_fd_pr__res_generic_m5_EGUVWD_0
timestamp 1696854327
transform 0 1 17009 1 0 48772
box -500 -257 500 257
use sky130_fd_pr__res_generic_m5_EGUVWD  sky130_fd_pr__res_generic_m5_EGUVWD_1
timestamp 1696854327
transform 0 1 17009 1 0 55228
box -500 -257 500 257
use sky130_fd_pr__res_generic_m5_EGUVWD  sky130_fd_pr__res_generic_m5_EGUVWD_2
timestamp 1696854327
transform 1 0 5927 0 -1 34243
box -500 -257 500 257
use sky130_fd_pr__res_generic_m5_EGUVWD  sky130_fd_pr__res_generic_m5_EGUVWD_3
timestamp 1696854327
transform 1 0 -5927 0 -1 34243
box -500 -257 500 257
<< labels >>
flabel metal5 17266 54728 17366 55728 0 FreeSans 1600 0 0 0 p1
port 1 nsew
flabel metal5 17266 48272 17366 49272 0 FreeSans 1600 0 0 0 p2
port 2 nsew
flabel metal5 5427 33886 6427 33986 0 FreeSans 1600 0 0 0 s1
port 3 nsew
flabel metal5 -6427 33886 -5427 33986 0 FreeSans 1600 0 0 0 s2
port 4 nsew
flabel metal5 16752 51500 16852 52500 0 FreeSans 1600 0 0 0 pm
port 5 nsew
<< end >>
