magic
tech sky130A
timestamp 1689171970
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 0.170 l 0.170 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 12.8 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
