magic
tech sky130A
timestamp 1694441024
<< error_p >>
rect -278 -144 -249 -141
rect 250 -144 279 -141
rect -278 -161 -272 -144
rect 250 -161 256 -144
rect -278 -164 -249 -161
rect 250 -164 279 -161
<< pwell >>
rect -371 -230 372 240
<< nmos >>
rect -271 -125 -256 125
rect -223 -125 -208 125
rect -175 -125 -160 125
rect -127 -125 -112 125
rect -79 -125 -64 125
rect -31 -125 -16 125
rect 17 -125 32 125
rect 65 -125 80 125
rect 113 -125 128 125
rect 161 -125 176 125
rect 209 -125 224 125
rect 257 -125 272 125
<< ndiff >>
rect -302 119 -271 125
rect -302 -119 -296 119
rect -279 -119 -271 119
rect -302 -125 -271 -119
rect -256 119 -223 125
rect -256 -119 -248 119
rect -231 -119 -223 119
rect -256 -125 -223 -119
rect -208 119 -175 125
rect -208 -119 -200 119
rect -183 -119 -175 119
rect -208 -125 -175 -119
rect -160 119 -127 125
rect -160 -119 -152 119
rect -135 -119 -127 119
rect -160 -125 -127 -119
rect -112 119 -79 125
rect -112 -119 -104 119
rect -87 -119 -79 119
rect -112 -125 -79 -119
rect -64 119 -31 125
rect -64 -119 -56 119
rect -39 -119 -31 119
rect -64 -125 -31 -119
rect -16 119 17 125
rect -16 -119 -8 119
rect 9 -119 17 119
rect -16 -125 17 -119
rect 32 119 65 125
rect 32 -119 40 119
rect 57 -119 65 119
rect 32 -125 65 -119
rect 80 119 113 125
rect 80 -119 88 119
rect 105 -119 113 119
rect 80 -125 113 -119
rect 128 119 161 125
rect 128 -119 136 119
rect 153 -119 161 119
rect 128 -125 161 -119
rect 176 119 209 125
rect 176 -119 184 119
rect 201 -119 209 119
rect 176 -125 209 -119
rect 224 119 257 125
rect 224 -119 232 119
rect 249 -119 257 119
rect 224 -125 257 -119
rect 272 119 303 125
rect 272 -119 280 119
rect 297 -119 303 119
rect 272 -125 303 -119
<< ndiffc >>
rect -296 -119 -279 119
rect -248 -119 -231 119
rect -200 -119 -183 119
rect -152 -119 -135 119
rect -104 -119 -87 119
rect -56 -119 -39 119
rect -8 -119 9 119
rect 40 -119 57 119
rect 88 -119 105 119
rect 136 -119 153 119
rect 184 -119 201 119
rect 232 -119 249 119
rect 280 -119 297 119
<< psubdiff >>
rect -353 195 -305 212
rect 306 195 354 212
rect -353 164 -336 195
rect 337 164 354 195
rect -353 -195 -336 -164
rect 337 -195 354 -164
rect -353 -212 -305 -195
rect 306 -212 354 -195
<< psubdiffcont >>
rect -305 195 306 212
rect -353 -164 -336 164
rect 337 -164 354 164
rect -305 -212 306 -195
<< poly >>
rect -271 125 -256 138
rect -223 125 -208 138
rect -175 125 -160 138
rect -127 125 -112 138
rect -79 125 -64 138
rect -31 125 -16 138
rect 17 125 32 138
rect 65 125 80 138
rect 113 125 128 138
rect 161 125 176 138
rect 209 125 224 138
rect 257 125 272 138
rect -271 -136 -256 -125
rect -223 -136 -208 -125
rect -175 -136 -160 -125
rect -280 -144 -247 -136
rect -280 -161 -272 -144
rect -255 -161 -247 -144
rect -280 -169 -247 -161
rect -223 -144 -160 -136
rect -223 -161 -215 -144
rect -168 -161 -160 -144
rect -223 -169 -160 -161
rect -127 -136 -112 -125
rect -79 -136 -64 -125
rect -127 -144 -64 -136
rect -127 -161 -119 -144
rect -72 -161 -64 -144
rect -127 -169 -64 -161
rect -31 -136 -16 -125
rect 17 -136 32 -125
rect -31 -144 32 -136
rect -31 -161 -23 -144
rect 24 -161 32 -144
rect -31 -169 32 -161
rect 65 -136 80 -125
rect 113 -136 128 -125
rect 65 -144 128 -136
rect 65 -161 73 -144
rect 120 -161 128 -144
rect 65 -169 128 -161
rect 161 -136 176 -125
rect 209 -136 224 -125
rect 257 -136 272 -125
rect 161 -144 224 -136
rect 161 -161 169 -144
rect 216 -161 224 -144
rect 161 -169 224 -161
rect 248 -144 281 -136
rect 248 -161 256 -144
rect 273 -161 281 -144
rect 248 -169 281 -161
<< polycont >>
rect -272 -161 -255 -144
rect -215 -161 -168 -144
rect -119 -161 -72 -144
rect -23 -161 24 -144
rect 73 -161 120 -144
rect 169 -161 216 -144
rect 256 -161 273 -144
<< locali >>
rect -353 195 -305 212
rect 306 195 354 212
rect -353 164 -336 195
rect 337 164 354 195
rect -296 119 -279 127
rect -296 -127 -279 -119
rect -248 119 -231 127
rect -248 -127 -231 -119
rect -200 119 -183 127
rect -200 -127 -183 -119
rect -152 119 -135 127
rect -152 -127 -135 -119
rect -104 119 -87 127
rect -104 -127 -87 -119
rect -56 119 -39 127
rect -56 -127 -39 -119
rect -8 119 9 127
rect -8 -127 9 -119
rect 40 119 57 127
rect 40 -127 57 -119
rect 88 119 105 127
rect 88 -127 105 -119
rect 136 119 153 127
rect 136 -127 153 -119
rect 184 119 201 127
rect 184 -127 201 -119
rect 232 119 249 127
rect 232 -127 249 -119
rect 280 119 297 127
rect 280 -127 297 -119
rect -280 -161 -272 -144
rect -255 -161 -247 -144
rect -223 -161 -215 -144
rect -168 -161 -160 -144
rect -127 -161 -119 -144
rect -72 -161 -64 -144
rect -31 -161 -23 -144
rect 24 -161 32 -144
rect 65 -161 73 -144
rect 120 -161 128 -144
rect 161 -161 169 -144
rect 216 -161 224 -144
rect 248 -161 256 -144
rect 273 -161 281 -144
rect -353 -195 -336 -164
rect 337 -195 354 -164
rect -353 -212 -305 -195
rect 306 -212 354 -195
<< viali >>
rect -296 -119 -279 119
rect -248 -119 -231 119
rect -200 -119 -183 119
rect -152 -119 -135 119
rect -104 -119 -87 119
rect -56 -119 -39 119
rect -8 -119 9 119
rect 40 -119 57 119
rect 88 -119 105 119
rect 136 -119 153 119
rect 184 -119 201 119
rect 232 -119 249 119
rect 280 -119 297 119
rect -272 -161 -255 -144
rect -215 -161 -168 -144
rect -119 -161 -72 -144
rect -23 -161 24 -144
rect 73 -161 120 -144
rect 169 -161 216 -144
rect 256 -161 273 -144
<< metal1 >>
rect -299 119 -276 125
rect -299 -119 -296 119
rect -279 -119 -276 119
rect -299 -125 -276 -119
rect -251 119 -228 125
rect -251 -119 -248 119
rect -231 -119 -228 119
rect -251 -125 -228 -119
rect -203 119 -180 125
rect -203 -119 -200 119
rect -183 -119 -180 119
rect -203 -125 -180 -119
rect -155 119 -132 125
rect -155 -119 -152 119
rect -135 -119 -132 119
rect -155 -125 -132 -119
rect -107 119 -84 125
rect -107 -119 -104 119
rect -87 -119 -84 119
rect -107 -125 -84 -119
rect -59 119 -36 125
rect -59 -119 -56 119
rect -39 -119 -36 119
rect -59 -125 -36 -119
rect -11 119 12 125
rect -11 -119 -8 119
rect 9 -119 12 119
rect -11 -125 12 -119
rect 37 119 60 125
rect 37 -119 40 119
rect 57 -119 60 119
rect 37 -125 60 -119
rect 85 119 108 125
rect 85 -119 88 119
rect 105 -119 108 119
rect 85 -125 108 -119
rect 133 119 156 125
rect 133 -119 136 119
rect 153 -119 156 119
rect 133 -125 156 -119
rect 181 119 204 125
rect 181 -119 184 119
rect 201 -119 204 119
rect 181 -125 204 -119
rect 229 119 252 125
rect 229 -119 232 119
rect 249 -119 252 119
rect 229 -125 252 -119
rect 277 119 300 125
rect 277 -119 280 119
rect 297 -119 300 119
rect 277 -125 300 -119
rect -278 -144 -249 -141
rect -278 -161 -272 -144
rect -255 -161 -249 -144
rect -278 -164 -249 -161
rect -221 -144 -162 -141
rect -221 -161 -215 -144
rect -168 -161 -162 -144
rect -221 -164 -162 -161
rect -125 -144 -66 -141
rect -125 -161 -119 -144
rect -72 -161 -66 -144
rect -125 -164 -66 -161
rect -29 -144 30 -141
rect -29 -161 -23 -144
rect 24 -161 30 -144
rect -29 -164 30 -161
rect 67 -144 126 -141
rect 67 -161 73 -144
rect 120 -161 126 -144
rect 67 -164 126 -161
rect 163 -144 222 -141
rect 163 -161 169 -144
rect 216 -161 222 -144
rect 163 -164 222 -161
rect 250 -144 279 -141
rect 250 -161 256 -144
rect 273 -161 279 -144
rect 250 -164 279 -161
<< properties >>
string FIXED_BBOX -345 -203 345 203
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
