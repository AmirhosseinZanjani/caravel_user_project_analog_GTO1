* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_564V44 a_n2867_n400# a_n1519_n497# a_n487_n497# a_n1261_n497#
+ a_487_n400# a_n29_n400# a_2609_n497# a_545_n497# a_2351_n497# a_2293_n400# a_n1835_n400#
+ a_1577_n497# a_n2809_n497# a_1519_n400# a_n803_n400# a_n2093_n400# a_n2551_n497#
+ a_1261_n400# a_n1777_n497# a_n1319_n400# a_29_n497# a_n287_n400# a_n1061_n400# a_n745_n497#
+ a_2809_n400# a_803_n497# a_n2035_n497# a_745_n400# a_2551_n400# a_1777_n400# a_n2609_n400#
+ a_1835_n497# a_n229_n497# a_n2351_n400# a_287_n497# a_n1003_n497# a_2093_n497# a_229_n400#
+ a_n1577_n400# a_2035_n400# a_n545_n400# a_1319_n497# w_n3005_n619# a_n2293_n497#
+ a_1061_n497# a_1003_n400#
X0 a_n1577_n400# a_n1777_n497# a_n1835_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_1519_n400# a_1319_n497# a_1261_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n1061_n400# a_n1261_n497# a_n1319_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_745_n400# a_545_n497# a_487_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_1003_n400# a_803_n497# a_745_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_487_n400# a_287_n497# a_229_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_1777_n400# a_1577_n497# a_1519_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_2035_n400# a_1835_n497# a_1777_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n2609_n400# a_n2809_n497# a_n2867_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X9 a_1261_n400# a_1061_n497# a_1003_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n1835_n400# a_n2035_n497# a_n2093_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_2809_n400# a_2609_n497# a_2551_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X12 a_n2351_n400# a_n2551_n497# a_n2609_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_n2093_n400# a_n2293_n497# a_n2351_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_n29_n400# a_n229_n497# a_n287_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_229_n400# a_29_n497# a_n29_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_n1319_n400# a_n1519_n497# a_n1577_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_2551_n400# a_2351_n497# a_2293_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_n545_n400# a_n745_n497# a_n803_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_n287_n400# a_n487_n497# a_n545_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_2293_n400# a_2093_n497# a_2035_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_n803_n400# a_n1003_n497# a_n1061_n400# w_n3005_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_ACGK3H a_n2093_n200# a_1261_n200# a_1319_n288# a_n2293_n288#
+ a_n1319_n200# a_1061_n288# a_n287_n200# a_n1061_n200# a_n1519_n288# a_2809_n200#
+ a_745_n200# a_n487_n288# a_n1261_n288# a_2551_n200# a_2609_n288# a_545_n288# a_1777_n200#
+ a_n2609_n200# a_2351_n288# a_n2351_n200# a_1577_n288# a_229_n200# a_n2809_n288#
+ a_n1577_n200# a_n2551_n288# a_2035_n200# a_n545_n200# a_29_n288# a_n1777_n288# a_n745_n288#
+ a_n2969_n374# a_1003_n200# a_803_n288# a_n2035_n288# a_n2867_n200# a_487_n200# a_n29_n200#
+ a_1835_n288# a_2293_n200# a_n229_n288# a_n1835_n200# a_287_n288# a_n1003_n288# a_n803_n200#
+ a_2093_n288# a_1519_n200#
X0 a_1003_n200# a_803_n288# a_745_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_745_n200# a_545_n288# a_487_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_487_n200# a_287_n288# a_229_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1777_n200# a_1577_n288# a_1519_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_2035_n200# a_1835_n288# a_1777_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n2609_n200# a_n2809_n288# a_n2867_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X6 a_1261_n200# a_1061_n288# a_1003_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n1835_n200# a_n2035_n288# a_n2093_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_2809_n200# a_2609_n288# a_2551_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X9 a_n2351_n200# a_n2551_n288# a_n2609_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n2093_n200# a_n2293_n288# a_n2351_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n29_n200# a_n229_n288# a_n287_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_229_n200# a_29_n288# a_n29_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_n1319_n200# a_n1519_n288# a_n1577_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_2551_n200# a_2351_n288# a_2293_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_n545_n200# a_n745_n288# a_n803_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_n287_n200# a_n487_n288# a_n545_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_2293_n200# a_2093_n288# a_2035_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_n803_n200# a_n1003_n288# a_n1061_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_n1577_n200# a_n1777_n288# a_n1835_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_1519_n200# a_1319_n288# a_1261_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X21 a_n1061_n200# a_n1261_n288# a_n1319_n200# a_n2969_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt Quantizer Vss InP InN OP ON vdd Clk VSUBS
Xsky130_fd_pr__pfet_01v8_564V44_0 NodeA1 vdd Clk Clk vdd vdd vdd Clk Clk NodeA2 NodeA1
+ Clk vdd vdd ON vdd Clk OP Clk ON ON ON vdd Clk NodeA2 Clk Clk OP vdd NodeA2 vdd
+ Clk OP NodeA1 Clk Clk Clk OP vdd vdd vdd vdd vdd Clk Clk vdd sky130_fd_pr__pfet_01v8_564V44
Xsky130_fd_pr__nfet_01v8_ACGK3H_0 ON NodeA2 ON Vss NodeA1 InN Vss m1_1798_488# OP
+ Vss NodeA2 Clk InP OP Vss InN Vss ON Vss Vss Vss Vss Vss ON Vss OP m1_1798_488#
+ Clk Vss InP Vss m1_1798_488# InN Vss Vss m1_1798_488# m1_1798_488# Vss Vss Clk Vss
+ Clk InP NodeA1 Vss OP sky130_fd_pr__nfet_01v8_ACGK3H
.ends

.subckt sky130_fd_pr__pfet_01v8_T2K7LE a_10261_n3500# a_8203_n3500# a_8261_n3597#
+ a_n16493_n3500# a_12319_n3500# a_12377_n3597# a_n2029_n3597# a_n6203_n3500# a_n14377_n3597#
+ a_n10319_n3500# a_14435_n3597# a_29_n3597# a_n16435_n3597# a_2087_n3597# a_2029_n3500#
+ a_14377_n3500# a_n4087_n3597# a_n8261_n3500# a_4145_n3597# a_n12377_n3500# a_16435_n3500#
+ a_n6145_n3597# a_6203_n3597# a_n14435_n3500# a_10319_n3597# a_n10261_n3597# a_n8203_n3597#
+ w_n16631_n3719# a_n12319_n3597# a_4087_n3500# a_6145_n3500# a_n29_n3500# a_n2087_n3500#
+ a_n4145_n3500#
X0 a_14377_n3500# a_12377_n3597# a_12319_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X1 a_10261_n3500# a_8261_n3597# a_8203_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X2 a_n14435_n3500# a_n16435_n3597# a_n16493_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=10.15 ps=70.58 w=35 l=10
X3 a_4087_n3500# a_2087_n3597# a_2029_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X4 a_n6203_n3500# a_n8203_n3597# a_n8261_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X5 a_n29_n3500# a_n2029_n3597# a_n2087_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X6 a_2029_n3500# a_29_n3597# a_n29_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X7 a_16435_n3500# a_14435_n3597# a_14377_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=10.15 pd=70.58 as=5.075 ps=35.29 w=35 l=10
X8 a_n2087_n3500# a_n4087_n3597# a_n4145_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X9 a_6145_n3500# a_4145_n3597# a_4087_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X10 a_n10319_n3500# a_n12319_n3597# a_n12377_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X11 a_n12377_n3500# a_n14377_n3597# a_n14435_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X12 a_n8261_n3500# a_n10261_n3597# a_n10319_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X13 a_n4145_n3500# a_n6145_n3597# a_n6203_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X14 a_12319_n3500# a_10319_n3597# a_10261_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
X15 a_8203_n3500# a_6203_n3597# a_6145_n3500# w_n16631_n3719# sky130_fd_pr__pfet_01v8 ad=5.075 pd=35.29 as=5.075 ps=35.29 w=35 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_NJ4FLX a_n14377_n2088# a_n30841_n2088# a_14435_n2088#
+ a_29_n2088# a_28783_n2000# a_n14435_n2000# a_20551_n2000# a_n16435_n2088# a_4087_n2000#
+ a_n26783_n2000# a_26783_n2088# a_32899_n2000# a_22609_n2000# a_n33059_n2174# a_n28783_n2088#
+ a_n2087_n2000# a_2087_n2088# a_6145_n2000# a_n29_n2000# a_n20609_n2000# a_n28841_n2000#
+ a_n30899_n2000# a_30899_n2088# a_28841_n2088# a_20609_n2088# a_n20551_n2088# a_n4087_n2088#
+ a_18493_n2000# a_n22609_n2088# a_n32899_n2088# a_10261_n2000# a_n4145_n2000# a_4145_n2088#
+ a_8203_n2000# a_n32957_n2000# a_16493_n2088# a_n16493_n2000# a_n6145_n2088# a_12319_n2000#
+ a_n6203_n2000# a_6203_n2088# a_n18493_n2088# a_18551_n2088# a_10319_n2088# a_n10261_n2088#
+ a_24667_n2000# a_n10319_n2000# a_n18551_n2000# a_n8203_n2088# a_n12319_n2088# a_n22667_n2000#
+ a_22667_n2088# a_26725_n2000# a_n24667_n2088# a_2029_n2000# a_n24725_n2000# a_24725_n2088#
+ a_30841_n2000# a_14377_n2000# a_n26725_n2088# a_n8261_n2000# a_8261_n2088# a_12377_n2088#
+ a_16435_n2000# a_n12377_n2000# a_n2029_n2088#
X0 a_n26783_n2000# a_n28783_n2088# a_n28841_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X1 a_n6203_n2000# a_n8203_n2088# a_n8261_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X2 a_n29_n2000# a_n2029_n2088# a_n2087_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X3 a_2029_n2000# a_29_n2088# a_n29_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X4 a_16435_n2000# a_14435_n2088# a_14377_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X5 a_n2087_n2000# a_n4087_n2088# a_n4145_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X6 a_6145_n2000# a_4145_n2088# a_4087_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X7 a_n10319_n2000# a_n12319_n2088# a_n12377_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X8 a_18493_n2000# a_16493_n2088# a_16435_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X9 a_n30899_n2000# a_n32899_n2088# a_n32957_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=10
X10 a_n12377_n2000# a_n14377_n2088# a_n14435_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X11 a_26725_n2000# a_24725_n2088# a_24667_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X12 a_n20609_n2000# a_n22609_n2088# a_n22667_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X13 a_28783_n2000# a_26783_n2088# a_26725_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X14 a_n22667_n2000# a_n24667_n2088# a_n24725_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X15 a_n8261_n2000# a_n10261_n2088# a_n10319_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X16 a_n4145_n2000# a_n6145_n2088# a_n6203_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X17 a_12319_n2000# a_10319_n2088# a_10261_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X18 a_8203_n2000# a_6203_n2088# a_6145_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X19 a_32899_n2000# a_30899_n2088# a_30841_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=10
X20 a_20551_n2000# a_18551_n2088# a_18493_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X21 a_14377_n2000# a_12377_n2088# a_12319_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X22 a_n18551_n2000# a_n20551_n2088# a_n20609_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X23 a_10261_n2000# a_8261_n2088# a_8203_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X24 a_n14435_n2000# a_n16435_n2088# a_n16493_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X25 a_4087_n2000# a_2087_n2088# a_2029_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X26 a_22609_n2000# a_20609_n2088# a_20551_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X27 a_n16493_n2000# a_n18493_n2088# a_n18551_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X28 a_30841_n2000# a_28841_n2088# a_28783_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X29 a_24667_n2000# a_22667_n2088# a_22609_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X30 a_n28841_n2000# a_n30841_n2088# a_n30899_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
X31 a_n24725_n2000# a_n26725_n2088# a_n26783_n2000# a_n33059_n2174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=10
.ends

.subckt integrator vdd BiasP1 InP InN OP ON BiasN1 BiasN2 BiasTail vss BiasP2 VSUBS
Xsky130_fd_pr__pfet_01v8_T2K7LE_0 NodeA vdd BiasP2 vdd ON BiasP1 BiasP2 NodeB BiasP1
+ NodeB vdd BiasP2 vdd BiasP2 NodeA NodeA BiasP2 vdd BiasP2 OP vdd BiasP2 BiasP2 NodeB
+ BiasP1 BiasP2 BiasP2 vdd BiasP1 vdd NodeA vdd NodeB vdd sky130_fd_pr__pfet_01v8_T2K7LE
Xsky130_fd_pr__nfet_01v8_NJ4FLX_0 InP BiasN1 InN ON vss Tail1 ON InP Tail1 m1_2132_284#
+ BiasN1 vss m1_55634_430# vss BiasN1 m1_26822_988# BiasTail m1_26822_988# vss OP
+ vss m1_2132_284# vss BiasN1 BiasN2 vss BiasTail vss BiasN2 vss Tail1 Tail1 BiasTail
+ vss vss vss NodeB BiasTail NodeA m1_26822_988# vss vss vss InN vss vss Tail1 vss
+ vss InP m1_2132_284# BiasN1 m1_55634_430# BiasN1 m1_26822_988# vss BiasN1 m1_55634_430#
+ Tail1 BiasN1 vss vss InN NodeA NodeB OP sky130_fd_pr__nfet_01v8_NJ4FLX
X0 ON OP sky130_fd_pr__cap_mim_m3_2 l=14.62 w=31.83
X1 OP ON sky130_fd_pr__cap_mim_m3_2 l=14.62 w=31.83
.ends

.subckt merg1b integrator_0/InN integrator_0/BiasP2 Quantizer_0/vdd Quantizer_0/InP
+ Quantizer_0/Vss Quantizer_0/InN Quantizer_0/Clk integrator_0/InP integrator_0/BiasN1
+ Quantizer_0/ON integrator_0/BiasN2 Quantizer_0/OP integrator_0/BiasP1
XQuantizer_0 Quantizer_0/Vss Quantizer_0/InP Quantizer_0/InN Quantizer_0/OP Quantizer_0/ON
+ Quantizer_0/vdd Quantizer_0/Clk VSUBS Quantizer
Xintegrator_0 Quantizer_0/vdd integrator_0/BiasP1 integrator_0/InP integrator_0/InN
+ Quantizer_0/OP Quantizer_0/ON integrator_0/BiasN1 integrator_0/BiasN2 integrator_0/BiasTail
+ Quantizer_0/Vss integrator_0/BiasP2 VSUBS integrator
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4524 pd=4.52 as=0.2262 ps=2.26 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4524 pd=4.52 as=0.2262 ps=2.26 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4524 pd=4.52 as=0.2262 ps=2.26 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR CLK D RESET_B Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4524 pd=4.52 as=0.2262 ps=2.26 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR X A1 S A0 VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=2
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=8
X2 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15 M=8
X3 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15 M=2
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15 M=4
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VGND VPWR VNB VPB
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 VGND LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__nor2b_2 VGND VPWR Y A B_N VNB VPB
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X4 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR A X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=16
X2 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15 M=4
X3 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15 M=16
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR X A B VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR CLK D RESET_B Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X11 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X15 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X16 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X17 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X22 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND X A VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=4
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR CLK D RESET_B Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15 M=4
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15 M=4
X11 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X15 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X16 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X17 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X22 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt adc_bridge VDD adc_cfg1[0] adc_cfg1[10] adc_cfg1[11] adc_cfg1[12] adc_cfg1[13]
+ adc_cfg1[14] adc_cfg1[15] adc_cfg1[1] adc_cfg1[2] adc_cfg1[3] adc_cfg1[4] adc_cfg1[5]
+ adc_cfg1[6] adc_cfg1[7] adc_cfg1[8] adc_cfg1[9] adc_cfg2[0] adc_cfg2[10] adc_cfg2[11]
+ adc_cfg2[12] adc_cfg2[13] adc_cfg2[14] adc_cfg2[15] adc_cfg2[1] adc_cfg2[2] adc_cfg2[3]
+ adc_cfg2[4] adc_cfg2[5] adc_cfg2[6] adc_cfg2[7] adc_cfg2[8] adc_cfg2[9] adc_conv_finished
+ adc_conv_finished_osr adc_res[0] adc_res[10] adc_res[11] adc_res[12] adc_res[13]
+ adc_res[14] adc_res[15] adc_res[1] adc_res[2] adc_res[3] adc_res[4] adc_res[5] adc_res[6]
+ adc_res[7] adc_res[8] adc_res[9] clk conv_finish dat_i dat_o load rst_n tie0 tie1
+ VSS
XFILLER_0_94_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_134_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Left_246 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_116_Left_255 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_432_ VSS VDD clknet_3_4_0_clk _076_ net63 adc_cfg_load_r\[23\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Left_264 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_363_ VSS VDD clknet_3_1_0_clk _027_ net58 net35 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_294_ VSS VDD _055_ _146_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_134_Left_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_89_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_89_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_129_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_125_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_346_ VSS VDD _081_ _172_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_415_ VSS VDD clknet_3_0_0_clk _059_ net58 adc_cfg_load_r\[6\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_277_ VSS VDD _138_ adc_cfg_load_r\[27\] _130_ net40 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_75_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_75_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_115_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_131_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_200_ VSS VDD _001_ _097_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_137_Right_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_20_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_136_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_45_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_329_ VSS VDD _164_ adc_cfg_load_r\[20\] net71 adc_cfg_load_r\[21\] VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_104_Right_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk clknet_3_1_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_56_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_21_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_97_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_34_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_26_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_107_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_128_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput42 VDD VSS adc_cfg2[13] net42 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput31 VDD VSS adc_cfg1[3] net31 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput53 VSS VDD net53 adc_cfg2[9] VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_23_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_362_ VSS VDD clknet_3_1_0_clk _026_ net58 net34 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_431_ VSS VDD clknet_3_4_0_clk _075_ net63 adc_cfg_load_r\[22\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_293_ VSS VDD _146_ adc_cfg_load_r\[2\] net70 adc_cfg_load_r\[3\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_64_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_104_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_118_Right_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_54_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_345_ VSS VDD _172_ adc_cfg_load_r\[28\] net72 adc_cfg_load_r\[29\] VSS VDD sky130_fd_sc_hd__mux2_1
X_414_ VSS VDD clknet_3_0_0_clk _058_ net58 adc_cfg_load_r\[5\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_276_ VSS VDD _046_ _137_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_40_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Right_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Right_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_136_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_61_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_259_ VSS VDD _038_ _128_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_328_ VSS VDD _072_ _163_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_101_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_19_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_31_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_72_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_122_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_137_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_137_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_27_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_26_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold20 net95 net52 VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_clk clknet_3_0_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xoutput43 VSS VDD net43 adc_cfg2[14] VSS VDD sky130_fd_sc_hd__clkbuf_4
Xoutput54 VSS VDD net54 conv_finish VSS VDD sky130_fd_sc_hd__clkbuf_4
Xoutput32 VDD VSS adc_cfg1[4] net32 VSS VDD sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Right_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_94_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Right_86 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_292_ VSS VDD _054_ _145_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_361_ VSS VDD clknet_3_1_0_clk _025_ net61 net33 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_430_ VSS VDD clknet_3_4_0_clk _074_ net62 adc_cfg_load_r\[21\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_95_Right_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_178 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Left_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_80_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_104_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_89_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_89_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_196 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_413_ VSS VDD clknet_3_0_0_clk _057_ net60 adc_cfg_load_r\[4\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_344_ VSS VDD _080_ _171_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_275_ VSS VDD _137_ adc_cfg_load_r\[26\] _130_ net39 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_59_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_115_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_65_Left_204 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_49_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_57_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Left_213 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Left_222 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_29_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Left_231 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_189_ VSS VDD _092_ net12 net67 net79 VSS VDD sky130_fd_sc_hd__mux2_1
X_258_ VSS VDD _128_ adc_cfg_load_r\[18\] _119_ net46 VSS VDD sky130_fd_sc_hd__mux2_1
X_327_ VSS VDD _163_ adc_cfg_load_r\[19\] net71 adc_cfg_load_r\[20\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_35_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_112_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_115_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_97_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_97_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_46_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold10 net85 adc_res_r\[13\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Left_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_6_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_67_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_107_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_16_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutput44 VDD VSS adc_cfg2[15] net44 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput55 VSS VDD net55 dat_o VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput22 VSS VDD net22 adc_cfg1[0] VSS VDD sky130_fd_sc_hd__clkbuf_4
Xoutput33 VDD VSS adc_cfg1[5] net33 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_78_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_78_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_94_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_134_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_7_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_291_ VSS VDD _145_ adc_cfg_load_r\[1\] net69 adc_cfg_load_r\[2\] VSS VDD sky130_fd_sc_hd__mux2_1
X_360_ VSS VDD clknet_3_1_0_clk _024_ net59 net32 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_103_Left_242 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_132_Right_132 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_120_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_13_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_13_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_89_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Left_251 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Left_260 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_412_ VSS VDD clknet_3_0_0_clk _056_ net59 adc_cfg_load_r\[3\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_343_ VSS VDD _171_ adc_cfg_load_r\[27\] net72 adc_cfg_load_r\[28\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_50_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_274_ VSS VDD _045_ _136_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_115_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_24_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_131_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_326_ VSS VDD _071_ _162_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_188_ VSS VDD _013_ _091_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_9_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_257_ VSS VDD _037_ _127_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_56_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_309_ VSS VDD _154_ adc_cfg_load_r\[10\] net72 adc_cfg_load_r\[11\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_21_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_108_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_97_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xhold11 net86 adc_res_r\[7\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_123_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_32_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput23 VDD VSS adc_cfg1[10] net23 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput34 VDD VSS adc_cfg1[6] net34 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput45 VDD VSS adc_cfg2[1] net45 VSS VDD sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_113_Right_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_53_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_118_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_94_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_290_ VSS VDD _053_ _144_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_13_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_129_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_411_ VSS VDD clknet_3_0_0_clk _055_ net59 adc_cfg_load_r\[2\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_342_ VSS VDD _079_ _170_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_273_ VSS VDD _136_ adc_cfg_load_r\[25\] _130_ net53 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_91_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_138_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_131_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_40_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_81_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_325_ VSS VDD _162_ adc_cfg_load_r\[18\] net71 adc_cfg_load_r\[19\] VSS VDD sky130_fd_sc_hd__mux2_1
X_187_ VSS VDD _091_ net11 net67 net84 VSS VDD sky130_fd_sc_hd__mux2_1
X_256_ VSS VDD _127_ adc_cfg_load_r\[17\] _119_ net45 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_126_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_19_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_51_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_62_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_56_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_72_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_308_ VSS VDD _062_ _153_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_239_ VSS VDD _118_ adc_cfg_load_r\[9\] _108_ net37 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_137_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_137_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Right_127 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold12 net87 adc_res_r\[11\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_107_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_107_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_16_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_120_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_25_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput24 VDD VSS adc_cfg1[11] net24 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput35 VDD VSS adc_cfg1[7] net35 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput46 VDD VSS adc_cfg2[2] net46 VSS VDD sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_134_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_27_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Right_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_134_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_46_Right_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Right_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_84_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Right_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_64_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_73_Right_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_82_Right_82 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_89_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_129_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_129_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_26_Left_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_92_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_44_Left_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_192 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_410_ VSS VDD clknet_3_0_0_clk _054_ net59 adc_cfg_load_r\[1\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_272_ VSS VDD _044_ _135_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_341_ VSS VDD _170_ adc_cfg_load_r\[26\] net72 adc_cfg_load_r\[27\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_59_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_115_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_115_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_24_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Left_200 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xfanout70 VSS VDD net20 net70 VSS VDD sky130_fd_sc_hd__clkbuf_4
X_255_ VSS VDD _036_ _126_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_324_ VSS VDD _070_ _161_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_108_Right_108 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_19_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_186_ VSS VDD _012_ _090_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_126_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_55_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_76_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_72_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_307_ VSS VDD _153_ adc_cfg_load_r\[9\] net72 adc_cfg_load_r\[10\] VSS VDD sky130_fd_sc_hd__mux2_1
X_238_ VSS VDD _028_ _117_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_137_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_46_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xhold13 net88 adc_res_r\[9\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_16_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_123_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_32_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_113_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput25 VDD VSS adc_cfg1[12] net25 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput36 VDD VSS adc_cfg1[8] net36 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput47 VDD VSS adc_cfg2[3] net47 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_78_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_27_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_134_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Left_238 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_7_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_80_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_13_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_104_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_85_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_271_ VSS VDD _135_ adc_cfg_load_r\[24\] _130_ net95 VSS VDD sky130_fd_sc_hd__mux2_1
X_340_ VSS VDD _078_ _169_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_24_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_131_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_40_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_185_ VSS VDD _090_ net10 net67 net82 VSS VDD sky130_fd_sc_hd__mux2_1
Xfanout60 VDD VSS net60 net21 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout71 VSS VDD net73 net71 VSS VDD sky130_fd_sc_hd__clkbuf_4
X_254_ VSS VDD _126_ adc_cfg_load_r\[16\] _119_ net38 VSS VDD sky130_fd_sc_hd__mux2_1
X_323_ VSS VDD _161_ adc_cfg_load_r\[17\] net71 adc_cfg_load_r\[18\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_101_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_86_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_126_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_35_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_48_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_306_ VSS VDD _061_ _152_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_237_ VSS VDD _117_ adc_cfg_load_r\[8\] _108_ net36 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_62_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Left_219 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_102_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_442__74 net74 _442__74/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xhold14 net89 adc_res_r\[14\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_119_Left_258 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_267 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_Left_276 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_83_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_32_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_106_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput26 VDD VSS adc_cfg1[13] net26 VSS VDD sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xoutput37 VSS VDD net37 adc_cfg1[9] VSS VDD sky130_fd_sc_hd__clkbuf_4
Xoutput48 VDD VSS adc_cfg2[4] net48 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_78_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_94_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_7_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_120_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_129_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_38_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_78_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_270_ VSS VDD _043_ _134_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_399_ VSS VDD clknet_3_3_0_clk _001_ net57 adc_res_r\[10\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_122_Right_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_322_ VSS VDD _069_ _160_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_100_Left_239 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_253_ VSS VDD _035_ _125_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_184_ VSS VDD _011_ _089_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xfanout61 VSS VDD net63 net61 VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout72 VSS VDD net73 net72 VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_86_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_136_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_51_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_51_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_305_ VSS VDD _152_ adc_cfg_load_r\[8\] net70 adc_cfg_load_r\[9\] VSS VDD sky130_fd_sc_hd__mux2_1
X_236_ VSS VDD _027_ _116_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_137_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_46_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_60_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold15 net90 adc_res_r\[17\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_219_ VSS VDD _107_ adc_cfg_written_r net71 VSS VDD sky130_fd_sc_hd__nor2b_2
XFILLER_0_57_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput27 VSS VDD net27 adc_cfg1[14] VSS VDD sky130_fd_sc_hd__clkbuf_4
Xoutput38 VDD VSS adc_cfg2[0] net38 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput49 VDD VSS adc_cfg2[5] net49 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_118_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_27_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_94_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_134_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk VSS VDD clk clknet_0_clk VSS VDD sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_15_Right_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Right_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Right_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_89_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_136_Right_136 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_129_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_38_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_54_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_60_Right_60 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_152 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_161 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_170 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_115_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_398_ VSS VDD clknet_3_3_0_clk _018_ net56 adc_res_r\[9\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_252_ VSS VDD _125_ adc_cfg_load_r\[15\] _119_ net28 VSS VDD sky130_fd_sc_hd__mux2_1
Xfanout73 VSS VDD net20 net73 VSS VDD sky130_fd_sc_hd__clkbuf_4
X_321_ VSS VDD _160_ adc_cfg_load_r\[16\] net71 adc_cfg_load_r\[17\] VSS VDD sky130_fd_sc_hd__mux2_1
Xfanout62 VSS VDD net63 net62 VSS VDD sky130_fd_sc_hd__clkbuf_4
X_183_ VSS VDD _089_ net3 net67 net91 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_126_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_35_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_129_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_235_ VSS VDD _116_ adc_cfg_load_r\[7\] _108_ net35 VSS VDD sky130_fd_sc_hd__mux2_1
X_304_ VSS VDD _060_ _151_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_46_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_62_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold16 net91 adc_res_r\[3\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_89_Right_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Right_98 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_144 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_123_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_16_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_218_ VSS VDD _019_ _106_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput28 VDD VSS adc_cfg1[15] net28 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput39 VSS VDD net39 adc_cfg2[10] VSS VDD sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_117_Right_117 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_134_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_111_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_7_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_68_Left_207 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_108_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Left_216 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Left_234 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_104_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_54_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_70_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_24_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_131_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_397_ VSS VDD clknet_3_3_0_clk _017_ net56 adc_res_r\[8\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_65_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_121_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_83_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_251_ VSS VDD _034_ _124_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_320_ VSS VDD _068_ _159_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_182_ VSS VDD _010_ _088_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xfanout63 VSS VDD net21 net63 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_51_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Left_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_92_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_112_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_234_ VSS VDD _026_ _115_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_303_ VSS VDD _151_ adc_cfg_load_r\[7\] net69 adc_cfg_load_r\[8\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_62_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold17 net92 adc_res_r\[18\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_106_Left_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_32_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_217_ VSS VDD _106_ net71 adc_cfg_written_r VSS VDD sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_115_Left_254 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_124_Left_263 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_73_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Left_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xoutput29 VDD VSS adc_cfg1[1] net29 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_68_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_104_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_104_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_120_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_129_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_54_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_396_ VSS VDD clknet_3_2_0_clk _016_ net56 adc_res_r\[7\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_49_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_49_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_4_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_81_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_76_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_250_ VSS VDD _124_ adc_cfg_load_r\[14\] _119_ net27 VSS VDD sky130_fd_sc_hd__mux2_1
Xfanout64 VSS VDD net66 net64 VSS VDD sky130_fd_sc_hd__clkbuf_4
X_181_ _088_ net67 net93 VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_0_19_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_379_ VSS VDD clknet_3_6_0_clk _043_ net62 net51 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_116_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_302_ VSS VDD _059_ _150_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_233_ VSS VDD _115_ adc_cfg_load_r\[6\] _108_ net34 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_137_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_46_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_134_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold18 net93 adc_res_r\[2\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_107_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_216_ VSS VDD _009_ _105_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_57_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_131_Right_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_118_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_84_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_120_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_38_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_79_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_21_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_115_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_395_ VSS VDD clknet_3_2_0_clk _015_ net56 adc_res_r\[6\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout65 VSS VDD net66 net65 VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_180_ VSS VDD _000_ _087_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_378_ VSS VDD clknet_3_6_0_clk _042_ net62 net50 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_132_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_301_ VSS VDD _150_ adc_cfg_load_r\[6\] net69 adc_cfg_load_r\[7\] VSS VDD sky130_fd_sc_hd__mux2_1
X_232_ VSS VDD _025_ _114_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_62_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_127_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Right_112 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_102_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Right_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_87_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold19 net94 adc_res_r\[16\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Right_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Right_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_123_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_215_ _105_ net69 net77 VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_85_Right_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_73_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Right_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_140 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_177 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_186 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Left_195 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_118_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_134_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_84_56 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_99_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_13_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_212 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_54_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Left_221 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_79_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Left_230 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_119_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_95_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_131_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_394_ VSS VDD clknet_3_2_0_clk _014_ net56 adc_res_r\[5\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_30_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_126_Right_126 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xfanout66 VDD VSS net66 net21 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_126_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_51_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_377_ VSS VDD clknet_3_6_0_clk _041_ net62 net49 VSS VDD sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_92_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_81_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_21_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_300_ VSS VDD _058_ _149_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_231_ VSS VDD _114_ adc_cfg_load_r\[5\] _108_ net33 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_62_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_429_ VSS VDD clknet_3_4_0_clk _073_ net62 adc_cfg_load_r\[20\] VSS VDD sky130_fd_sc_hd__dfrtp_1
Xinput1 VSS VDD net1 adc_conv_finished VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_214_ VSS VDD _008_ _104_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_44_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_102_Left_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_111_Left_250 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_134_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_17_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_129_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Right_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_79_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_102_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Right_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_28_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_135_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_24_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_393_ VSS VDD clknet_3_2_0_clk _013_ net56 adc_res_r\[4\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_49_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout56 VSS VDD net60 net56 VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout67 VSS VDD net70 net67 VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_376_ VSS VDD clknet_3_6_0_clk _040_ net62 net48 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_25_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_74_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_230_ VSS VDD _024_ _113_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_428_ VSS VDD clknet_3_4_0_clk _072_ net62 adc_cfg_load_r\[19\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_359_ VSS VDD clknet_3_1_0_clk _023_ net59 net31 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput2 VSS VDD net2 adc_conv_finished_osr VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_213_ VSS VDD _104_ net9 net69 net92 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_57_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_132_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_138_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_37_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_27_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_33_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_130_Left_269 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_110_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_110_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_95_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_392_ VSS VDD clknet_3_2_0_clk _012_ net56 adc_res_r\[3\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_65_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_105_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout68 VSS VDD net70 net68 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout57 VSS VDD net60 net57 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_375_ VSS VDD clknet_3_6_0_clk _039_ net62 net47 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_92_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_132_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_41_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_5_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_358_ VSS VDD clknet_3_1_0_clk _022_ net59 net30 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_427_ VSS VDD clknet_3_4_0_clk _071_ net63 adc_cfg_load_r\[18\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_289_ VSS VDD _144_ adc_cfg_load_r\[0\] net69 adc_cfg_load_r\[1\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_102_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Right_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xinput3 VSS VDD net3 adc_res[0] VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_212_ VSS VDD _007_ _103_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_45_Right_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_73_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_125_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_113_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Right_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_155 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_164 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_173 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_43_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Left_182 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_108_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Left_191 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_84_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_38_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_54_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_121_Right_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_119_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_69_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_97_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_391_ VSS VDD clknet_3_2_0_clk _011_ net56 adc_res_r\[2\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_81_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_39_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout69 VSS VDD net70 net69 VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout58 VSS VDD net60 net58 VSS VDD sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_8_Left_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_443_ VDD VSS tie1 net75 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_51_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_374_ VSS VDD clknet_3_6_0_clk _038_ net61 net46 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_92_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_46_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_62_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_11_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_357_ VSS VDD clknet_3_1_0_clk _021_ net59 net29 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_426_ VSS VDD clknet_3_4_0_clk _070_ net61 adc_cfg_load_r\[17\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_288_ VSS VDD _052_ _143_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput4 VSS VDD net4 adc_res[10] VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_89_Left_228 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Left_237 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_211_ VSS VDD _103_ net8 net69 net90 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_118_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_113_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_409_ VSS VDD clknet_3_1_0_clk _053_ net59 adc_cfg_load_r\[0\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_138_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Right_135 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_102_Right_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_108_56 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_42_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_54_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_70_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_119_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_28_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_390_ VSS VDD clknet_3_2_0_clk _010_ net56 adc_res_r\[1\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_71_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout59 VSS VDD net60 net59 VSS VDD sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_70_Left_209 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Left_248 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_442_ VDD VSS tie0 net74 VSS VDD sky130_fd_sc_hd__buf_2
X_373_ VSS VDD clknet_3_6_0_clk _037_ net61 net45 VSS VDD sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_118_Left_257 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_132_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Left_266 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_25_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_136_Left_275 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_66_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_82_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_356_ VSS VDD clknet_3_0_0_clk _020_ net59 net22 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_287_ VSS VDD _143_ adc_cfg_load_r\[32\] _107_ conv_finish_sel VSS VDD sky130_fd_sc_hd__mux2_1
X_425_ VSS VDD clknet_3_4_0_clk _069_ net61 adc_cfg_load_r\[16\] VSS VDD sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_116_Right_116 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_87_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_127_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput5 VSS VDD net5 adc_res[11] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_72_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_210_ VSS VDD _006_ _102_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_113_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_22_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_408_ VSS VDD clknet_3_0_0_clk net69 net58 adc_res_r\[19\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_339_ VSS VDD _169_ adc_cfg_load_r\[25\] net72 adc_cfg_load_r\[26\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_138_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_47_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_68_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_17_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_130_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_33_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_35_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_70_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_95_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_65_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_121_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_121_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_441_ VSS VDD clknet_3_4_0_clk _085_ net61 adc_cfg_load_r\[32\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_372_ VSS VDD clknet_3_6_0_clk _036_ net61 net38 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_25_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_132_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_41_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_424_ VSS VDD clknet_3_5_0_clk _068_ net66 adc_cfg_load_r\[15\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_286_ VSS VDD _051_ _142_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_355_ VSS VDD clknet_3_4_0_clk _019_ net61 adc_cfg_written_r VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput6 VSS VDD net6 adc_res[12] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_73_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_22_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Right_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_407_ VSS VDD clknet_3_1_0_clk _009_ net58 adc_res_r\[18\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_338_ VSS VDD _077_ _168_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_269_ VSS VDD _134_ adc_cfg_load_r\[23\] _130_ net51 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_138_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Right_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_50_Right_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_68_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_84_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_160 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_33_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_123_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput20 VSS VDD load net20 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_99_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_119_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_28_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Right_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_81_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_39_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_95_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_371_ VSS VDD clknet_3_7_0_clk _035_ net65 net28 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_440_ VSS VDD clknet_3_4_0_clk _084_ net61 adc_cfg_load_r\[31\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_79_Right_79 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Right_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_76_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_92_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_97_Right_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_143 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_41_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_10_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Left_198 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Right_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_423_ VSS VDD clknet_3_5_0_clk _067_ net66 adc_cfg_load_r\[14\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_354_ VSS VDD _085_ _176_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_285_ VSS VDD _142_ adc_cfg_load_r\[31\] _107_ net44 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_36_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_127_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput7 VSS VDD net7 adc_res[13] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_206 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_215 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Left_224 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_406_ VSS VDD clknet_3_1_0_clk _008_ net58 adc_res_r\[17\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_337_ VSS VDD _168_ adc_cfg_load_r\[24\] net72 adc_cfg_load_r\[25\] VSS VDD sky130_fd_sc_hd__mux2_1
X_199_ VSS VDD _097_ net17 net68 net87 VSS VDD sky130_fd_sc_hd__mux2_1
X_268_ VSS VDD _042_ _133_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_94_Left_233 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_138_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_17_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_84_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput21 VSS VDD rst_n net21 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_0_116_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput10 VSS VDD net10 adc_res[1] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_119_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_28_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_44_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_8_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_179 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_105_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_39_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_111_Right_111 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_88_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_370_ VSS VDD clknet_3_7_0_clk _034_ net65 net27 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_25_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_92_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_132_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_66_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_105_Left_244 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_114_Left_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Left_262 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_132_Left_271 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_422_ VSS VDD clknet_3_5_0_clk _066_ net66 adc_cfg_load_r\[13\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_284_ VSS VDD _050_ _141_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_353_ VSS VDD _176_ adc_cfg_load_r\[32\] net71 net19 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_87_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_36_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput8 VSS VDD net8 adc_res[14] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_113_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_405_ VSS VDD clknet_3_1_0_clk _007_ net58 adc_res_r\[16\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_267_ VSS VDD _133_ adc_cfg_load_r\[22\] _130_ net50 VSS VDD sky130_fd_sc_hd__mux2_1
X_336_ VSS VDD _076_ _167_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_198_ VSS VDD _018_ _096_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_138_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_33_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_319_ VSS VDD _159_ adc_cfg_load_r\[15\] net73 adc_cfg_load_r\[16\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_109_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput11 VSS VDD net11 adc_res[2] VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_125_Right_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_95_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_60_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_109_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_33_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_121_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_55_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_96_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_25_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_132_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_41_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_421_ VSS VDD clknet_3_5_0_clk _065_ net65 adc_cfg_load_r\[12\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_283_ VSS VDD _141_ adc_cfg_load_r\[30\] _107_ net43 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_11_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_352_ VSS VDD _084_ _175_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_127_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput9 VSS VDD net9 adc_res[15] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_404_ VSS VDD clknet_3_3_0_clk _006_ net57 adc_res_r\[15\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_197_ VSS VDD _096_ net16 net67 net80 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_22_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_266_ VSS VDD _041_ _132_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_335_ VSS VDD _167_ adc_cfg_load_r\[23\] net73 adc_cfg_load_r\[24\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_98_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_63_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_106_Right_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_318_ VSS VDD _067_ _158_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_249_ VSS VDD _033_ _123_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput12 VSS VDD net12 adc_res[3] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_110_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_119_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_121_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_39_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold1 net76 adc_res_r\[1\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_71_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Right_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_66_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Right_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_167 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_93_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Right_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_176 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_420_ VSS VDD clknet_3_5_0_clk _064_ net65 adc_cfg_load_r\[11\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_351_ VSS VDD _175_ adc_cfg_load_r\[31\] net71 adc_cfg_load_r\[32\] VSS VDD sky130_fd_sc_hd__mux2_1
X_282_ VSS VDD _049_ _140_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_46_Left_185 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_102_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_127_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_194 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_403_ VSS VDD clknet_3_3_0_clk _005_ net57 adc_res_r\[14\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_334_ VSS VDD _075_ _166_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_196_ VSS VDD _017_ _095_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_265_ VSS VDD _132_ adc_cfg_load_r\[21\] _130_ net49 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_138_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Left_202 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_211 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_81_Left_220 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_108_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_317_ VSS VDD _158_ adc_cfg_load_r\[14\] net73 adc_cfg_load_r\[15\] VSS VDD sky130_fd_sc_hd__mux2_1
Xinput13 VSS VDD net13 adc_res[4] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_248_ VSS VDD _123_ adc_cfg_load_r\[13\] _119_ net26 VSS VDD sky130_fd_sc_hd__mux2_1
X_179_ VSS VDD _087_ net67 net76 VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_0_74_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_90_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_110_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_28_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_114_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_69_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_19_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_105_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold2 net77 adc_res_r\[19\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_116_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_82_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_350_ VSS VDD _083_ _174_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_281_ VSS VDD _140_ adc_cfg_load_r\[29\] _130_ net42 VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_101_Left_240 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_36_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_77_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_113_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_402_ VSS VDD clknet_3_3_0_clk _004_ net57 adc_res_r\[13\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_264_ VSS VDD _040_ _131_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_333_ VSS VDD _166_ adc_cfg_load_r\[22\] net73 adc_cfg_load_r\[23\] VSS VDD sky130_fd_sc_hd__mux2_1
X_195_ VSS VDD _095_ net15 net67 net88 VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_120_Right_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_49_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_108_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_316_ VSS VDD _066_ _157_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_247_ VSS VDD _032_ _122_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput14 VSS VDD net14 adc_res[5] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_178_ VSS VDD _086_ net54 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_0_90_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_107_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_8_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_69_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_85_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_109_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_121_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold3 net78 adc_res_r\[15\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_116_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_132_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_41_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_79_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_134_Right_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_280_ VSS VDD _048_ _139_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_52_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_101_Right_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_77_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_93_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_401_ VSS VDD clknet_3_3_0_clk _003_ net57 adc_res_r\[12\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_263_ VSS VDD _131_ adc_cfg_load_r\[20\] _130_ net48 VSS VDD sky130_fd_sc_hd__mux2_1
X_332_ VSS VDD _074_ _165_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_194_ VSS VDD _016_ _094_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_88_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Left_259 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_124_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_315_ VSS VDD _157_ adc_cfg_load_r\[13\] net73 adc_cfg_load_r\[14\] VSS VDD sky130_fd_sc_hd__mux2_1
X_246_ VSS VDD _122_ adc_cfg_load_r\[12\] _119_ net25 VSS VDD sky130_fd_sc_hd__mux2_1
Xinput15 VSS VDD net15 adc_res[6] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_177_ VSS VDD _086_ net1 conv_finish_sel net2 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_61_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_119_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_8_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_229_ VSS VDD _113_ adc_cfg_load_r\[4\] _108_ net32 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_69_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold4 net79 adc_res_r\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_71_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_115_Right_115 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_111_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_96_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_136_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_24_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Right_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_132_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Right_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_106_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Right_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Right_62 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_154 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_127_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_163 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_172 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_77_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Left_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_133_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Left_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_400_ VSS VDD clknet_3_3_0_clk _002_ net57 adc_res_r\[11\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_331_ VSS VDD _165_ adc_cfg_load_r\[21\] net71 adc_cfg_load_r\[22\] VSS VDD sky130_fd_sc_hd__mux2_1
X_262_ VSS VDD _107_ _130_ VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_193_ VSS VDD _094_ net14 net67 net81 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_138_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_17_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_314_ VSS VDD _065_ _156_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_245_ VSS VDD _031_ _121_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput16 VSS VDD net16 adc_res[7] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_114_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_23_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_99_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_54_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Right_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_28_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_135_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_146 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_228_ VSS VDD _023_ _112_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_85_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_85_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_30_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold5 net80 adc_res_r\[10\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_112_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_111_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_17_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_79_Left_218 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_25_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_88_Left_227 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Left_236 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_36_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_77_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_84_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_6_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_330_ VSS VDD _073_ _164_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_192_ VSS VDD _015_ _093_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_261_ VSS VDD _039_ _129_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_12_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_103_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_313_ VSS VDD _156_ adc_cfg_load_r\[12\] net73 adc_cfg_load_r\[13\] VSS VDD sky130_fd_sc_hd__mux2_1
X_244_ VSS VDD _121_ adc_cfg_load_r\[11\] _119_ net24 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_33_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput17 VSS VDD net17 adc_res[8] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_3_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_47_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_64_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_28_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_44_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_227_ VSS VDD _112_ adc_cfg_load_r\[3\] _108_ net31 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_109_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_108_Left_247 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Left_256 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Left_265 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Left_274 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xhold6 net81 adc_res_r\[8\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_111_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_20_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_105_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_29_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_96_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_41_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_82_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_106_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_36_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_52_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_77_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_260_ VSS VDD _129_ adc_cfg_load_r\[19\] _119_ net47 VSS VDD sky130_fd_sc_hd__mux2_1
X_191_ VSS VDD _093_ net13 net67 net86 VSS VDD sky130_fd_sc_hd__mux2_1
X_389_ VSS VDD clknet_3_2_0_clk _000_ net56 net55 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_312_ VSS VDD _064_ _155_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_243_ VSS VDD _030_ _120_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput18 VSS VDD net18 adc_res[9] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_114_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_90_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_99_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_110_Right_110 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_44_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_8_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_60_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_226_ VSS VDD _022_ _111_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_109_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_39_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xhold7 net82 adc_res_r\[4\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
X_209_ VSS VDD _102_ net7 net69 net94 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_136_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_15_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_122_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_56_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_72_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_40_Right_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_52_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_77_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_117_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_26_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_190_ VSS VDD _014_ _092_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_Right_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_12_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_388_ VSS VDD clknet_3_6_0_clk _052_ net61 conv_finish_sel VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_311_ VSS VDD _155_ adc_cfg_load_r\[11\] net72 adc_cfg_load_r\[12\] VSS VDD sky130_fd_sc_hd__mux2_1
X_242_ VSS VDD _120_ adc_cfg_load_r\[10\] _119_ net23 VSS VDD sky130_fd_sc_hd__mux2_1
Xinput19 VDD VSS net19 dat_i VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_58_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_114_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_23_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_130_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_60_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Right_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_225_ VSS VDD _111_ adc_cfg_load_r\[2\] _108_ net30 VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_78_Right_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_85_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_125_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_109_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_87_Right_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Right_96 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_52_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Left_188 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xhold8 net83 adc_res_r\[12\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_111_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_111_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_20_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_208_ VSS VDD _005_ _101_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Left_205 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_15_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_110_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_31_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Left_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Left_223 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Right_138 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_232 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Right_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_93_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_42_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_clk clknet_3_7_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_63_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_387_ VSS VDD clknet_3_7_0_clk _051_ net64 net44 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_128_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_82_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_310_ VSS VDD _063_ _154_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_30_Left_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_241_ VDD VSS _119_ _107_ VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_0_58_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_74_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_439_ VSS VDD clknet_3_5_0_clk _083_ net66 adc_cfg_load_r\[30\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_224_ VSS VDD _021_ _110_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_109_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_109_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_59_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_104_Left_243 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xhold9 net84 adc_res_r\[5\] VSS VDD VSS VDD sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_113_Left_252 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_71_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_122_Left_261 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_207_ VSS VDD _101_ net6 net68 net78 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_20_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_29_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_136_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_136_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_131_Left_270 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Right_119 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_66_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_82_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_106_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_31_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_103_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_117_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_26_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_67_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_386_ VSS VDD clknet_3_7_0_clk _050_ net64 net43 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_75_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_240_ VSS VDD _029_ _118_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_clk clknet_3_6_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_369_ VSS VDD clknet_3_7_0_clk _033_ net65 net26 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_438_ VSS VDD clknet_3_5_0_clk _082_ net66 adc_cfg_load_r\[29\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_223_ VSS VDD _110_ adc_cfg_load_r\[1\] _108_ net29 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_69_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_125_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_34_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_59_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_206_ VSS VDD _004_ _100_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_136_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_86_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_82_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_106_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_15_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_56_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_77_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_26_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_42_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_6_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_20_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_385_ VSS VDD clknet_3_7_0_clk _049_ net64 net42 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_88_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_37_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_53_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_114_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_23_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_90_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_368_ VSS VDD clknet_3_7_0_clk _032_ net65 net25 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_437_ VSS VDD clknet_3_5_0_clk _081_ net64 adc_cfg_load_r\[28\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_299_ VSS VDD _149_ adc_cfg_load_r\[5\] net69 adc_cfg_load_r\[6\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_104_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Right_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_222_ VSS VDD _020_ _109_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_47_Right_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_34_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_50_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Right_56 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Right_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_91_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_74_Right_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_clk clknet_3_5_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_18_Left_157 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_166 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_111_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_205_ VSS VDD _100_ net5 net68 net89 VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_36_Left_175 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_96_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Left_184 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_9_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_61_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_100_Right_100 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_50_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_122_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_31_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_201 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_98_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Left_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_93_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_117_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_42_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_6_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_13_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_384_ VSS VDD clknet_3_7_0_clk _048_ net64 net41 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_88_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_53_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_436_ VSS VDD clknet_3_5_0_clk _080_ net64 adc_cfg_load_r\[27\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_367_ VSS VDD clknet_3_7_0_clk _031_ net65 net24 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_298_ VSS VDD _057_ _148_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_80_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_114_Right_114 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_221_ VSS VDD _109_ adc_cfg_load_r\[0\] _108_ net22 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_100_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_109_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_419_ VSS VDD clknet_3_5_0_clk _063_ net65 adc_cfg_load_r\[10\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_119_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_204_ VSS VDD _003_ _099_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_96_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_29_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_136_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_61_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Left_139 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_56_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_clk clknet_3_4_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
X_443__75 _443__75/LO net75 VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_0_97_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_117_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_1 adc_cfg_load_r\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_101_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_383_ VSS VDD clknet_3_7_0_clk _047_ net64 net40 VSS VDD sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_128_Right_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_128_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_37_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_90_Left_229 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_129_Left_268 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_Left_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_366_ VSS VDD clknet_3_7_0_clk _030_ net65 net23 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_435_ VSS VDD clknet_3_7_0_clk _079_ net64 adc_cfg_load_r\[26\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_297_ VSS VDD _148_ adc_cfg_load_r\[4\] net70 adc_cfg_load_r\[5\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_64_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_64_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_220_ VSS VDD _107_ _108_ VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_18_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_125_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_418_ VSS VDD clknet_3_5_0_clk _062_ net65 adc_cfg_load_r\[9\] VSS VDD sky130_fd_sc_hd__dfrtp_4
X_349_ VSS VDD _174_ adc_cfg_load_r\[30\] net72 adc_cfg_load_r\[31\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_59_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_75_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_75_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_203_ VSS VDD _099_ net4 net68 net85 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_136_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_45_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_36_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_106_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_56_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_72_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_110_Left_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Right_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_26_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_133_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_2 net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_6_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_67_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_123_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_103_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_382_ VSS VDD clknet_3_7_0_clk _046_ net64 net39 VSS VDD sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_3_0_clk clknet_3_3_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
Xoutput50 VDD VSS adc_cfg2[6] net50 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_53_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_114_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_23_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_365_ VSS VDD clknet_3_1_0_clk _029_ net59 net37 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_296_ VSS VDD _056_ _147_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_434_ VSS VDD clknet_3_6_0_clk _078_ net64 adc_cfg_load_r\[25\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_80_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_66_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Right_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_348_ VSS VDD _082_ _173_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_279_ VSS VDD _139_ adc_cfg_load_r\[28\] _130_ net41 VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Right_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_417_ VSS VDD clknet_3_0_0_clk _061_ net60 adc_cfg_load_r\[8\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Right_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_91_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Right_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_111_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_202_ VSS VDD _002_ _098_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_61_Right_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_61_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_124_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Left_162 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Left_171 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_180 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_122_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_106_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_72_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Right_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_42_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_6_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_3 net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_83_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_96_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_381_ VSS VDD clknet_3_6_0_clk _045_ net62 net53 VSS VDD sky130_fd_sc_hd__dfrtp_1
Xoutput40 VDD VSS adc_cfg2[11] net40 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput51 VDD VSS adc_cfg2[7] net51 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_78_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Right_99 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_94_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_114_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_433_ VSS VDD clknet_3_4_0_clk _077_ net63 adc_cfg_load_r\[24\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_364_ VSS VDD clknet_3_1_0_clk _028_ net58 net36 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_295_ VSS VDD _147_ adc_cfg_load_r\[3\] net70 adc_cfg_load_r\[4\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_3_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_59_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_clk clknet_3_2_0_clk clknet_0_clk VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Left_208 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_416_ VSS VDD clknet_3_0_0_clk _060_ net58 adc_cfg_load_r\[7\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_347_ VSS VDD _173_ adc_cfg_load_r\[29\] net72 adc_cfg_load_r\[30\] VSS VDD sky130_fd_sc_hd__mux2_1
X_278_ VSS VDD _047_ _138_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Left_217 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_59_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_59_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_87_Left_226 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_91_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Left_235 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_201_ VSS VDD _098_ net18 net68 net83 VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_0_29_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_117_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_86_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_122_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_123_Right_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_97_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_41_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_117_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_67_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_67_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_60_Left_199 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_89_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_12_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_380_ VSS VDD clknet_3_6_0_clk _044_ net62 net52 VSS VDD sky130_fd_sc_hd__dfrtp_1
Xoutput41 VDD VSS adc_cfg2[12] net41 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput30 VDD VSS adc_cfg1[2] net30 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput52 VSS VDD net52 adc_cfg2[8] VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_37_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_78_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_94_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
.ends

.subckt sky130_fd_sc_hd__xor2_1 VPWR VGND A X B VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND A1 A2 X B1 B2 C1 VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND Y A VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15 M=2
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR A Y B VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR A B Y VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_2 VGND VPWR B1 B2 A2 A1 X C1 VNB VPB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3875 ps=1.775 w=1 l=0.15
X4 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X6 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.165 ps=1.33 w=1 l=0.15
X7 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3875 pd=1.775 as=0.1125 ps=1.225 w=1 l=0.15
X8 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X10 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23725 ps=2.03 w=0.65 l=0.15
X11 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR B Y A VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VGND VPWR A_N B Y VNB VPB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4524 pd=4.52 as=0.2262 ps=2.26 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 VGND VPWR X A2 A1 B1 C1 VNB VPB
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.13325 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.199875 pd=1.265 as=0.091 ps=0.93 w=0.65 l=0.15 M=2
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.199875 ps=1.265 w=0.65 l=0.15
X9 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_2 VPWR VGND A Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15 M=2
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=3
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR X A3 A2 A1 B1 B2 VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND B C A X VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR X A3 A2 A1 B1 VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VGND VPWR A B Y C VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X A B VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND A2 A1 B1 Y VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VGND VPWR A2 A1 Y B1 VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15 M=2
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=2
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15 M=2
X7 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND A X VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=6
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15 M=2
X2 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=6
X3 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR A X B_N VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR B1 B2 A2 A1 X C1 VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VGND VPWR A2 A1 B1 X VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15 M=2
X1 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15 M=2
X2 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X3 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X4 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X6 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VGND VPWR Y A B VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X C B A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_4 VPWR VGND A2 X A1 C1 B1 B2 VNB VPB
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15 M=2
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=4
X7 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X8 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X9 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
X10 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15 M=2
X11 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__nor3_1 VGND VPWR C B A Y VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR A1 A2 B1 X VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 VGND VPWR A Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt pfet_01v8_w500_l500_nf2 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26#
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND X A VNB VPB
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 nmoscap_top nmoscap_bot pwell sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
.ends

.subckt nfet_01v8_w500_l500_nf2 a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76# SUB a_129_n50#
X0 a_129_n50# a_29_n76# a_n29_n50# SUB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_n50# a_n129_n76# a_n187_n50# SUB sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt adc_vcm_generator clk phi2 phi1_n phi1 phi2_n vcm VDD mimtop1 mimtop2 mimbot1
+ VSS
Xsky130_fd_sc_hd__inv_1_4 VSS VDD clk sky130_fd_sc_hd__inv_1_4/Y VSS VDD sky130_fd_sc_hd__inv_1
Xpfet_01v8_w500_l500_nf2_0 mimtop2 vcm phi1_n VDD vcm phi1_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_1 mimtop1 vcm phi1_n VDD vcm phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_0 VDD VSS phi1 sky130_fd_sc_hd__inv_1_2/A VSS VDD sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_2 mimtop2 mimbot1 phi2_n VDD mimbot1 phi2_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_1 VDD VSS phi1_n sky130_fd_sc_hd__inv_1_2/Y VSS VDD sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_3 VDD mimtop1 phi2_n VDD mimtop1 phi2_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_4 mimbot1 VSS phi1_n VDD VSS phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_2 VDD VSS phi2 sky130_fd_sc_hd__inv_1_3/A VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_3 VDD VSS phi2_n sky130_fd_sc_hd__inv_1_3/Y VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__nand2_1_0/Y
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__nand2_1_1/Y
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 VDD VSS sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_3/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__dlymetal6s6s_1_4/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 VDD VSS sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|0] vcm VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|0] vcm VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|0] vcm VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|0] vcm VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|0] vcm VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|0] vcm VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|1] vcm VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|1] vcm VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|1] vcm VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|1] vcm VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|1] vcm VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|1] vcm VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|2] vcm VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|2] vcm VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|2] vcm VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|2] vcm VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|2] vcm VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|2] vcm VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|3] vcm VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|3] vcm VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|3] vcm VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|3] vcm VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|3] vcm VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|3] vcm VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|4] vcm VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|4] vcm VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|4] vcm VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|4] vcm VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|4] vcm VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|4] vcm VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top VSS
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xnfet_01v8_w500_l500_nf2_0 phi1 mimtop2 vcm phi1 VSS vcm nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_1 phi1 mimtop1 vcm phi1 VSS vcm nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_0 VSS VDD clk sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_2 phi2 mimtop2 mimbot1 phi2 VSS mimbot1 nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_3 phi2 VDD mimtop1 phi2 VSS mimtop1 nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_1 VSS VDD sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__nand2_1_1/Y
+ sky130_fd_sc_hd__inv_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_4 phi1 mimbot1 VSS phi1 VSS VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__inv_1_0 VSS VDD sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 VSS VDD sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_3/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 VSS VDD sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 VSS VDD sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15 M=2
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15 M=2
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15 M=2
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15 M=2
X4 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=2
X5 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND B1 A1 A2 X B2 VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND B D C A X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR A1 A2 Y B2 C1 B1 VNB VPB
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1652 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VGND VPWR C A Y B VNB VPB
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X4 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X5 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND A2 A1 B1 X VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 VGND VPWR X D C B A VNB VPB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinvlp_2 VGND VPWR A Y VNB VPB
X0 Y A a_150_67# VNB sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.67 as=0.066 ps=0.79 w=0.55 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.14 ps=1.28 w=1 l=0.25 M=2
X2 a_150_67# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.79 as=0.15675 ps=1.67 w=0.55 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR B C_N A X VNB VPB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VGND VPWR Y B C A_N VNB VPB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 VPWR VGND B1_N A2 Y A1 VNB VPB
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183125 ps=1.24 w=0.65 l=0.15 M=2
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=2
X5 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.06825 ps=0.86 w=0.65 l=0.15
X8 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183125 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X9 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VGND VPWR X A2 A1 B1_N VNB VPB
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR B2 A2 A1 B1 X VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 VGND VPWR Y B A VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=4
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15 M=4
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
.ends

.subckt sky130_fd_sc_hd__a221oi_1 VGND VPWR Y B1 C1 A1 A2 B2 VNB VPB
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.069875 pd=0.865 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.099125 ps=0.955 w=0.65 l=0.15
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.069875 ps=0.865 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.1525 ps=1.305 w=1 l=0.15
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 VPWR VGND A Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=6
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1659 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15 M=4
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt adc_array_matrix_12bit row_n[0] row_n[1] row_n[2] row_n[3] row_n[4] row_n[5]
+ row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12] row_n[13] row_n[14]
+ row_n[15] rowon_n[0] rowon_n[1] rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6]
+ rowon_n[7] rowon_n[8] rowon_n[9] rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13]
+ rowon_n[14] rowon_n[15] rowoff_n[0] rowoff_n[1] rowoff_n[2] rowoff_n[3] rowoff_n[4]
+ rowoff_n[5] rowoff_n[6] rowoff_n[7] rowoff_n[8] rowoff_n[9] rowoff_n[10] rowoff_n[11]
+ rowoff_n[12] rowoff_n[13] rowoff_n[14] rowoff_n[15] vcm sample sample_n col_n[31]
+ col_n[30] col_n[29] col_n[28] col_n[27] col_n[26] col_n[25] col_n[24] col_n[23]
+ col_n[22] col_n[21] col_n[20] col_n[19] col_n[18] col_n[17] col_n[16] col_n[15]
+ col_n[14] col_n[13] col_n[12] col_n[11] col_n[10] col_n[9] col_n[8] col_n[7] col_n[6]
+ col_n[5] col_n[4] col_n[3] col_n[2] col_n[1] col_n[0] en_bit_n[2] en_bit_n[1] en_bit_n[0]
+ en_C0_n sw sw_n analog_in col[0] col[1] col[2] col[3] col[4] col[5] col[6] col[7]
+ col[8] col[9] col[10] col[11] col[12] col[13] col[14] col[15] col[16] col[17] col[18]
+ col[19] col[20] col[21] col[22] col[23] col[24] col[25] col[26] col[27] col[28]
+ col[29] col[30] col[31] ctop VSS VDD
X0 a_3970_15182# a_2475_15206# a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1 a_3878_9158# a_2275_9182# a_3970_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2 VDD rowon_n[5] a_18938_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3 a_30986_7150# row_n[5] a_31478_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4 vcm a_2275_18218# a_32082_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_12002_2130# a_2475_2154# a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6 a_5374_4500# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X7 a_14410_15544# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X8 a_10906_12170# row_n[10] a_11398_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X9 a_35398_9198# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_17422_7512# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X11 a_18026_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X12 VSS row_n[4] a_9294_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_4370_15544# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X14 a_23046_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X15 a_22346_10202# rowon_n[8] a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X16 a_14922_11166# row_n[9] a_15414_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X17 a_15414_2492# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X18 a_4882_11166# row_n[9] a_5374_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X19 a_34394_2170# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_27062_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X21 VSS row_n[6] a_26362_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1957_14202# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X23 a_34090_3134# a_2475_3158# a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X24 a_1957_4162# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X25 a_26058_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X26 a_21342_2170# rowon_n[0] a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X27 a_35002_9158# row_n[7] a_35494_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X28 a_23350_18234# VDD a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X29 VSS row_n[13] a_20338_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_26970_14178# a_2275_14202# a_27062_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X31 a_11302_8194# rowon_n[6] a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X32 a_29982_4138# a_2275_4162# a_30074_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X33 a_12306_4178# rowon_n[2] a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X34 vcm a_2275_2154# a_13006_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 VDD rowon_n[3] a_22954_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X36 VSS row_n[12] a_24354_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_21342_11206# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_34394_10202# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_24962_17190# a_2275_17214# a_25054_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X40 a_18938_7150# a_2275_7174# a_19030_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X41 a_4274_13214# rowon_n[11] a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X42 a_14314_13214# rowon_n[11] a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X43 VSS row_n[8] a_11302_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_20034_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X45 a_21038_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X46 a_19430_18556# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X47 a_19030_14178# a_2475_14202# a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X48 a_11910_11166# a_2275_11190# a_12002_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X49 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X50 VDD rowon_n[14] a_22954_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X51 a_28978_14178# row_n[12] a_29470_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X52 a_20434_13536# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X53 a_33486_12532# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X54 vcm a_2275_10186# a_29070_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_20338_6186# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_15926_12170# a_2275_12194# a_16018_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X57 a_3270_7190# rowon_n[5] a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X58 VSS row_n[4] a_30378_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_4274_3174# rowon_n[1] a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X60 VDD rowon_n[2] a_11910_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X61 a_5886_12170# a_2275_12194# a_5978_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X62 VDD rowon_n[10] a_9902_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X63 a_16322_6186# rowon_n[4] a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X64 vcm a_2275_6170# a_24050_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_35398_18234# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15 M=2
X66 VDD rowon_n[9] a_3878_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X67 VDD rowon_n[9] a_13918_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X68 VDD rowon_n[4] a_5886_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X69 VSS VDD a_12306_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_30074_17190# a_2475_17214# a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X71 a_16018_7150# a_2475_7174# a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X72 a_26058_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X73 a_25054_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X74 a_13310_14218# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 VDD en_C0_n a_3878_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X76 a_30986_17190# row_n[15] a_31478_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X77 a_12002_16186# a_2475_16210# a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X78 a_34090_16186# a_2475_16210# a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X79 a_3270_14218# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X80 vcm a_2275_13198# a_31078_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_25358_4178# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X82 a_35002_16186# row_n[14] a_35494_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X83 a_10906_8154# row_n[6] a_11398_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X84 VSS row_n[6] a_34394_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X85 a_8290_5182# rowon_n[3] a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X86 a_9294_1166# VSS a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X87 VSS row_n[2] a_35398_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X88 a_9994_9158# a_2475_9182# a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X89 a_12402_16548# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X90 a_19334_16226# rowon_n[14] a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X91 a_20338_11206# rowon_n[9] a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X92 vcm a_2275_8178# a_28066_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 vcm a_2275_4162# a_29070_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X94 VSS a_2161_13198# a_2275_13198# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X95 a_25358_7190# rowon_n[5] a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X96 a_25054_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X97 a_13310_7190# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X98 a_29070_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X99 a_14314_3174# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X100 a_16018_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X101 a_33998_9158# a_2275_9182# a_34090_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X102 VDD rowon_n[1] a_7894_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X103 a_24962_4138# row_n[2] a_25454_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X104 a_5978_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X105 a_2874_7150# row_n[5] a_3366_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X106 vcm a_2275_7174# a_17022_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X107 a_35494_4500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X108 a_19942_11166# a_2275_11190# a_20034_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X109 a_32994_10162# a_2275_10186# a_33086_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X110 a_15926_6146# row_n[4] a_16418_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X111 a_34394_18234# VDD a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X112 a_27366_17230# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X113 VSS row_n[13] a_31382_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X114 a_13918_1126# VDD a_14410_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X115 VSS row_n[12] a_35398_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X116 a_32386_11206# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X117 a_6282_2170# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X118 a_22954_18194# a_2275_18218# a_23046_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X119 a_12306_14218# rowon_n[12] a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X120 a_18330_5182# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X121 a_19334_1166# en_bit_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15 M=2
X122 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X123 VDD rowon_n[15] a_29982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X124 a_26058_15182# a_2475_15206# a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X125 VSS en_bit_n[0] a_20338_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15 M=2
X126 vcm a_2275_11190# a_27062_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X127 a_7894_5142# row_n[3] a_8386_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X128 a_30378_1166# VSS a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X129 VDD rowon_n[14] a_33998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X130 a_26970_15182# row_n[13] a_27462_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X131 a_31478_13536# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X132 a_3878_13174# a_2275_13198# a_3970_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X133 a_13918_13174# a_2275_13198# a_14010_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X134 a_23046_5142# a_2475_5166# a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X135 VDD rowon_n[6] a_30986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X136 a_17934_3134# row_n[1] a_18426_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X137 a_29374_9198# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X138 a_29982_12170# row_n[10] a_30474_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X139 VSS row_n[1] a_24354_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X140 a_10394_7512# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X141 a_33390_7190# rowon_n[5] a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X142 a_34394_3174# rowon_n[1] a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X143 a_18330_11206# rowon_n[9] a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X144 a_10998_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X145 VSS row_n[7] a_14314_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X146 a_27062_7150# a_2475_7174# a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X147 a_28066_3134# a_2475_3158# a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X148 vcm a_2275_9182# a_32082_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X149 a_18938_18194# VDD a_19430_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X150 vcm a_2275_14202# a_8990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X151 vcm a_2275_14202# a_19030_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X152 a_4974_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X153 a_28978_9158# row_n[7] a_29470_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X154 a_8898_18194# VDD a_9390_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X155 a_22954_8154# a_2275_8178# a_23046_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X156 a_24450_1488# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X157 a_19030_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X158 VSS row_n[0] a_13310_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X159 a_23958_4138# a_2275_4162# a_24050_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X160 a_33086_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X161 a_23046_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X162 VSS VDD a_29374_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X163 a_14410_9520# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X164 a_15414_5504# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X165 VSS row_n[13] a_29374_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X166 a_33390_13214# rowon_n[11] a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X167 a_26362_12210# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X168 VSS row_n[8] a_30378_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X169 a_16018_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X170 VSS row_n[2] a_7286_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X171 a_30986_11166# a_2275_11190# a_31078_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X172 a_11910_7150# a_2275_7174# a_12002_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X173 VDD rowon_n[15] a_27974_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X174 a_25454_14540# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X175 a_35002_12170# a_2275_12194# a_35094_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X176 a_25054_10162# a_2475_10186# a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X177 a_27974_6146# a_2275_6170# a_28066_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X178 a_32082_1126# a_2475_1150# a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X179 a_5886_9158# a_2275_9182# a_5978_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X180 a_33998_18194# a_2275_18218# a_34090_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X181 a_29470_13536# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X182 VDD rowon_n[9] a_32994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X183 a_25966_10162# row_n[8] a_26458_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X184 a_32994_7150# row_n[5] a_33486_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X185 a_7382_4500# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X186 a_14010_2130# a_2475_2154# a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X187 a_30986_2130# row_n[0] a_31478_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X188 VDD rowon_n[0] a_18938_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X189 a_11910_14178# a_2275_14202# a_12002_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X190 VDD rowon_n[10] a_8898_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X191 a_16930_5142# a_2275_5166# a_17022_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X192 a_17422_2492# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X193 vcm a_2275_15206# a_23046_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X194 VSS row_n[6] a_28370_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X195 a_17022_17190# a_2475_17214# a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X196 a_8290_15222# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X197 a_18330_15222# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X198 a_6982_17190# a_2475_17214# a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X199 a_9902_17190# a_2275_17214# a_9994_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X200 a_1957_8178# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X201 a_23350_2170# rowon_n[0] a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X202 vcm a_2275_10186# a_14010_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X203 a_2966_9158# a_2475_9182# a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X204 a_2161_6170# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X205 a_7382_17552# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X206 a_17422_17552# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X207 a_3878_14178# row_n[12] a_4370_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X208 a_13918_14178# row_n[12] a_14410_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X209 a_25358_12210# rowon_n[10] a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X210 vcm a_2275_10186# a_3970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X211 a_13310_8194# rowon_n[6] a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X212 vcm a_2275_8178# a_21038_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X213 vcm a_2275_4162# a_22042_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X214 a_14314_4178# rowon_n[2] a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X215 a_17934_13174# row_n[11] a_18426_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X216 a_29374_11206# rowon_n[9] a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X217 a_31078_8154# a_2475_8178# a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X218 vcm a_2275_2154# a_15014_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_7894_13174# row_n[11] a_8386_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X220 VDD rowon_n[6] a_2874_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X221 a_23046_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X222 a_22042_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X223 VDD rowon_n[8] a_24962_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X224 VDD rowon_n[2] a_13918_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X225 vcm a_2275_18218# a_4974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X226 vcm a_2275_18218# a_15014_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X227 VSS row_n[15] a_23350_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X228 VSS row_n[4] a_32386_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X229 a_6282_3174# rowon_n[1] a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X230 vcm a_2275_6170# a_26058_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X231 VSS row_n[14] a_27366_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X232 a_31382_14218# rowon_n[12] a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X233 a_24354_13214# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X234 vcm a_2275_9182# a_3970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X235 VDD rowon_n[4] a_7894_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X236 a_2475_4162# a_1957_4162# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X237 a_32082_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X238 a_17326_15222# rowon_n[13] a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X239 a_11302_5182# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X240 a_12306_1166# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X241 a_28066_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X242 a_7286_15222# rowon_n[13] a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X243 a_19942_14178# a_2275_14202# a_20034_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X244 a_32994_13174# a_2275_13198# a_33086_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X245 a_18026_7150# a_2475_7174# a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X246 a_27062_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X247 VDD VDD a_25966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X248 a_3970_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X249 a_14010_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X250 a_23446_15544# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X251 VSS row_n[9] a_8290_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X252 VSS row_n[9] a_18330_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X253 a_23046_11166# a_2475_11190# a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X254 VDD VSS a_5886_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X255 a_23958_11166# row_n[9] a_24450_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X256 a_12914_8154# row_n[6] a_13406_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X257 VDD rowon_n[6] a_24962_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X258 VDD rowon_n[11] a_6890_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X259 VDD rowon_n[11] a_16930_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X260 a_10906_3134# row_n[1] a_11398_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X261 a_12306_17230# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X262 a_22346_9198# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X263 a_27366_7190# rowon_n[5] a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X264 a_16322_3174# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X265 vcm a_2275_4162# a_30074_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X266 a_16322_16226# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X267 vcm a_2275_16210# a_21038_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X268 a_15318_7190# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X269 a_15014_18194# a_2475_18218# a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X270 a_6282_16226# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X271 vcm a_2275_15206# a_34090_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X272 a_4882_7150# row_n[5] a_5374_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X273 a_4974_18194# a_2475_18218# a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X274 vcm a_2275_7174# a_19030_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X275 a_17934_6146# row_n[4] a_18426_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X276 a_21038_3134# a_2475_3158# a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X277 a_15414_18556# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X278 a_11910_15182# row_n[13] a_12402_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X279 vcm a_2275_11190# a_12002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X280 a_20034_7150# a_2475_7174# a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X281 a_2874_2130# row_n[0] a_3366_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X282 a_5374_18556# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X283 a_21950_9158# row_n[7] a_22442_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X284 a_15926_1126# VDD a_16418_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X285 a_8290_2170# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X286 a_28066_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X287 a_9902_2130# a_2275_2154# a_9994_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X288 VSS row_n[10] a_22346_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X289 VSS VDD a_22346_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X290 a_32386_1166# VSS a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X291 a_31382_5182# rowon_n[3] a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X292 a_26058_1126# a_2475_1150# a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X293 VSS VDD a_21342_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X294 a_25054_5142# a_2475_5166# a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X295 VDD rowon_n[12] a_20946_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X296 a_22346_14218# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X297 a_16322_10202# rowon_n[8] a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X298 VDD rowon_n[6] a_32994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X299 a_26970_7150# row_n[5] a_27462_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X300 a_6282_10202# rowon_n[8] a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X301 a_30074_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X302 a_22442_10524# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X303 a_20946_6146# a_2275_6170# a_21038_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X304 a_5278_16226# rowon_n[14] a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X305 a_15318_16226# rowon_n[14] a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X306 a_31078_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X307 VDD rowon_n[1] a_30986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X308 a_20338_17230# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X309 a_21438_16548# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X310 a_30986_14178# a_2275_14202# a_31078_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X311 a_18330_9198# rowon_n[7] a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X312 a_30378_9198# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X313 a_12402_7512# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X314 a_13006_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X315 VSS row_n[4] a_4274_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X316 a_6890_15182# a_2275_15206# a_6982_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X317 a_16930_15182# a_2275_15206# a_17022_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X318 vcm a_2275_9182# a_34090_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X319 a_29070_7150# a_2475_7174# a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X320 a_10394_2492# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X321 VSS row_n[13] a_4274_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X322 VSS row_n[13] a_14314_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X323 a_11302_12210# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X324 a_19942_15182# row_n[13] a_20434_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X325 a_15318_11206# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X326 vcm a_2275_11190# a_20034_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X327 a_6982_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X328 VSS row_n[6] a_21342_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X329 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X330 a_32994_14178# row_n[12] a_33486_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X331 a_14010_13174# a_2475_13198# a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X332 a_5278_11206# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X333 vcm a_2275_10186# a_33086_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X334 a_24962_8154# a_2275_8178# a_25054_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X335 VSS row_n[0] a_15318_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X336 a_25966_4138# a_2275_4162# a_26058_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X337 a_3970_13174# a_2475_13198# a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X338 VDD rowon_n[7] a_17934_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X339 a_29982_9158# row_n[7] a_30474_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X340 a_35094_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X341 VDD rowon_n[3] a_18938_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X342 a_30986_5142# row_n[3] a_31478_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X343 VDD rowon_n[15] a_2874_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X344 VDD rowon_n[15] a_12914_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X345 vcm a_2275_16210# a_32082_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X346 a_10394_14540# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X347 a_5978_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X348 a_14410_13536# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X349 a_10906_10162# row_n[8] a_11398_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X350 a_17422_5504# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X351 a_18026_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X352 VSS row_n[2] a_9294_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X353 a_4370_13536# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X354 VDD a_2161_7174# a_2275_7174# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X355 a_13918_7150# a_2275_7174# a_14010_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X356 VSS row_n[4] a_26362_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X357 a_1957_2154# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X358 a_26058_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X359 a_7894_9158# a_2275_9182# a_7986_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X360 a_35002_7150# row_n[5] a_35494_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X361 a_9390_4500# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X362 VSS VDD a_19334_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X363 a_23350_16226# rowon_n[14] a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X364 VSS row_n[11] a_20338_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X365 a_11302_6186# rowon_n[4] a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X366 VSS row_n[10] a_33390_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X367 a_32994_2130# row_n[0] a_33486_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X368 a_6890_2130# a_2275_2154# a_6982_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X369 a_10298_12210# rowon_n[10] a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X370 a_24962_15182# a_2275_15206# a_25054_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X371 a_18938_5142# a_2275_5166# a_19030_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X372 a_28066_12170# a_2475_12194# a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X373 a_4274_11206# rowon_n[9] a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X374 a_14314_11206# rowon_n[9] a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X375 a_10998_7150# a_2475_7174# a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X376 a_21038_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X377 a_20034_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X378 a_8990_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X379 a_19430_16548# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X380 VDD rowon_n[12] a_31990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X381 a_28978_12170# row_n[10] a_29470_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X382 a_20434_11528# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X383 a_33486_10524# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X384 a_20338_4178# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X385 a_3270_5182# rowon_n[3] a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X386 a_4274_1166# en_C0_n a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X387 VSS row_n[2] a_30378_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X388 a_31382_17230# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X389 VDD rowon_n[8] a_9902_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X390 a_4974_9158# a_2475_9182# a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X391 a_19030_2130# a_2475_2154# a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X392 a_16322_4178# rowon_n[2] a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X393 vcm a_2275_8178# a_23046_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X394 vcm a_2275_4162# a_24050_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X395 a_35398_16226# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X396 a_33086_8154# a_2475_8178# a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X397 VSS row_n[14] a_12306_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X398 a_20338_7190# rowon_n[5] a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X399 vcm a_2275_17214# a_26058_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X400 a_30074_15182# a_2475_15206# a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X401 a_24050_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X402 a_16018_5142# a_2475_5166# a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X403 a_25054_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X404 a_34090_14178# a_2475_14202# a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X405 VDD rowon_n[1] a_2874_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X406 a_19942_4138# row_n[2] a_20434_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X407 a_34490_18556# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X408 a_30986_15182# row_n[13] a_31478_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X409 a_12002_14178# a_2475_14202# a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X410 vcm a_2275_11190# a_31078_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X411 vcm a_2275_7174# a_12002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X412 a_30474_4500# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X413 VDD VDD a_10906_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X414 vcm a_2275_12194# a_17022_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X415 a_10906_6146# row_n[4] a_11398_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X416 VSS row_n[4] a_34394_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X417 a_8290_3174# rowon_n[1] a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X418 VDD rowon_n[2] a_15926_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X419 vcm a_2275_12194# a_6982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X420 a_19334_14218# rowon_n[12] a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X421 vcm a_2275_6170# a_28066_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X422 vcm a_2275_9182# a_5978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X423 a_21038_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X424 a_2475_8178# a_1957_8178# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X425 a_25358_5182# rowon_n[3] a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X426 a_13310_5182# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X427 a_14314_1166# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X428 a_29070_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X429 VDD VSS a_7894_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X430 VDD rowon_n[6] a_26970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X431 a_2874_5142# row_n[3] a_3366_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X432 vcm a_2275_5166# a_17022_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X433 a_30378_17230# rowon_n[15] a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X434 a_14922_8154# row_n[6] a_15414_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X435 a_3970_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X436 a_14010_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X437 a_34394_16226# rowon_n[14] a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X438 a_27366_15222# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X439 VSS row_n[11] a_31382_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X440 VDD rowon_n[1] a_24962_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X441 a_12914_3134# row_n[1] a_13406_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X442 a_24354_9198# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X443 VSS row_n[5] a_19334_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X444 a_29374_7190# rowon_n[5] a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X445 a_22954_16186# a_2275_16210# a_23046_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X446 a_18330_3174# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X447 a_6982_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X448 a_17022_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X449 a_26458_17552# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X450 VDD rowon_n[13] a_29982_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X451 a_26058_13174# a_2475_13198# a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X452 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X453 a_30378_12210# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X454 a_26970_13174# row_n[11] a_27462_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X455 a_31478_11528# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X456 a_22042_7150# a_2475_7174# a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X457 a_23046_3134# a_2475_3158# a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X458 VDD rowon_n[4] a_30986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X459 a_4882_2130# row_n[0] a_5374_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X460 vcm a_2275_12194# a_25054_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X461 a_23958_9158# row_n[7] a_24450_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X462 a_17934_1126# en_bit_n[1] a_18426_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X463 a_19334_18234# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X464 vcm a_2275_18218# a_24050_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X465 a_29982_10162# row_n[8] a_30474_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X466 a_9294_18234# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X467 VSS VDD a_24354_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X468 a_9390_14540# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X469 a_10394_5504# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X470 a_33390_5182# rowon_n[3] a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X471 a_28066_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X472 a_10998_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X473 a_28066_1126# a_2475_1150# a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X474 a_27062_5142# a_2475_5166# a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X475 a_19030_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X476 a_18938_16186# row_n[14] a_19430_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X477 a_28978_7150# row_n[5] a_29470_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X478 a_8898_16186# row_n[14] a_9390_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X479 a_22954_6146# a_2275_6170# a_23046_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X480 a_33086_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X481 a_26970_2130# row_n[0] a_27462_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X482 VDD rowon_n[1] a_32994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X483 a_28370_17230# rowon_n[15] a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X484 a_14410_7512# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X485 VSS row_n[11] a_29374_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X486 a_33390_11206# rowon_n[9] a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X487 a_26362_10202# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X488 a_15014_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X489 VSS a_2161_1150# a_2275_1150# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X490 a_16018_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X491 a_11910_5142# a_2275_5166# a_12002_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X492 a_12402_2492# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X493 a_9294_12210# rowon_n[10] a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X494 a_16930_10162# a_2275_10186# a_17022_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X495 a_8990_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X496 VSS row_n[6] a_23350_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X497 a_31382_2170# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X498 a_19334_2170# rowon_n[0] a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X499 VDD rowon_n[13] a_27974_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X500 a_25454_12532# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X501 a_6890_10162# a_2275_10186# a_6982_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X502 VSS row_n[0] a_17326_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X503 a_27974_4138# a_2275_4162# a_28066_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X504 a_33998_16186# a_2275_16210# a_34090_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X505 a_29470_11528# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X506 a_32994_5142# row_n[3] a_33486_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X507 a_7986_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X508 VDD rowon_n[8] a_8898_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X509 vcm a_2275_2154# a_9994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X510 VSS row_n[15] a_7286_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X511 VSS row_n[15] a_17326_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X512 a_22042_17190# a_2475_17214# a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X513 a_15926_7150# a_2275_7174# a_16018_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X514 a_16930_3134# a_2275_3158# a_17022_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X515 a_18330_13214# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X516 vcm a_2275_13198# a_23046_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X517 VSS row_n[4] a_28370_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X518 a_22954_17190# row_n[15] a_23446_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X519 a_17022_15182# a_2475_15206# a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X520 a_8290_13214# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X521 VSS row_n[7] a_6282_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X522 a_6982_15182# a_2475_15206# a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X523 a_9902_15182# a_2275_15206# a_9994_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X524 a_1957_6170# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X525 a_17422_15544# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X526 a_2161_4162# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X527 a_7382_15544# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X528 a_3878_12170# row_n[10] a_4370_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X529 a_13918_12170# row_n[10] a_14410_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X530 a_26058_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X531 a_25358_10202# rowon_n[8] a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X532 a_13310_6186# rowon_n[4] a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X533 vcm a_2275_6170# a_21038_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X534 a_17934_11166# row_n[9] a_18426_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X535 a_31078_6146# a_2475_6170# a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X536 a_35002_2130# row_n[0] a_35494_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X537 a_8898_2130# a_2275_2154# a_8990_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X538 a_7894_11166# row_n[9] a_8386_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X539 VDD rowon_n[4] a_2874_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X540 a_6378_9520# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X541 a_23046_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X542 a_13006_7150# a_2475_7174# a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X543 a_22042_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X544 vcm a_2275_17214# a_10998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X545 a_24962_10162# a_2275_10186# a_25054_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X546 VDD rowon_n[6] a_19942_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X547 a_26362_18234# VDD a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X548 vcm a_2275_16210# a_4974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X549 vcm a_2275_16210# a_15014_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X550 VSS row_n[13] a_23350_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X551 a_6982_9158# a_2475_9182# a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X552 a_6282_1166# VSS a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X553 VSS row_n[2] a_32386_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X554 vcm a_2275_8178# a_25054_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X555 vcm a_2275_4162# a_26058_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X556 VSS row_n[12] a_27366_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X557 a_24354_11206# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X558 a_35094_8154# a_2475_8178# a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X559 a_27974_17190# a_2275_17214# a_28066_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X560 a_5978_2130# a_2475_2154# a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X561 a_2475_2154# a_1957_2154# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X562 VDD rowon_n[15] a_21950_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X563 a_32082_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X564 a_17326_13214# rowon_n[11] a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X565 a_22346_7190# rowon_n[5] a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X566 a_11302_3174# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X567 a_7286_13214# rowon_n[11] a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X568 a_30986_9158# a_2275_9182# a_31078_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X569 a_10298_7190# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X570 a_18026_5142# a_2475_5166# a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X571 a_27062_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X572 VDD rowon_n[14] a_25966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X573 a_3970_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X574 a_14010_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X575 a_23446_13536# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X576 a_32482_4500# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X577 a_18938_12170# a_2275_12194# a_19030_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X578 vcm a_2275_7174# a_14010_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X579 a_12914_6146# row_n[4] a_13406_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X580 VDD rowon_n[4] a_24962_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X581 a_8898_12170# a_2275_12194# a_8990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X582 VDD rowon_n[9] a_6890_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X583 VDD rowon_n[9] a_16930_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X584 a_10906_1126# VDD a_11398_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X585 VSS VDD a_15318_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X586 a_20034_18194# a_2475_18218# a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X587 a_12306_15222# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X588 vcm a_2275_9182# a_7986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X589 a_3270_2170# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X590 VSS VDD a_5278_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X591 a_10998_17190# a_2475_17214# a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X592 a_33086_17190# a_2475_17214# a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X593 a_16322_1166# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X594 a_27366_5182# rowon_n[3] a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X595 a_20946_18194# VDD a_21438_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X596 a_16322_14218# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X597 vcm a_2275_14202# a_21038_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X598 a_5278_8194# rowon_n[6] a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X599 a_15318_5182# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X600 a_33998_17190# row_n[15] a_34490_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X601 a_15014_16186# a_2475_16210# a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X602 a_6282_14218# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X603 vcm a_2275_13198# a_34090_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X604 a_19430_8516# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X605 a_4882_5142# row_n[3] a_5374_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X606 vcm a_2275_2154# a_6982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X607 a_11398_17552# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X608 a_4974_16186# a_2475_16210# a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X609 VDD rowon_n[6] a_28978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X610 vcm a_2275_5166# a_19030_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X611 a_21038_1126# a_2475_1150# a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X612 a_20034_5142# a_2475_5166# a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X613 a_15414_16548# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X614 a_11910_13174# row_n[11] a_12402_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X615 VDD rowon_n[1] a_26970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X616 a_5374_16548# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X617 a_21950_7150# row_n[5] a_22442_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X618 a_14922_3134# row_n[1] a_15414_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X619 a_2475_16210# a_1957_16210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X620 a_28066_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X621 vcm a_2275_12194# a_9994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X622 a_26362_9198# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 VSS row_n[8] a_22346_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X624 a_22954_11166# a_2275_11190# a_23046_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X625 a_31382_3174# rowon_n[1] a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X626 a_25054_3134# a_2475_3158# a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X627 VSS row_n[14] a_21342_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X628 a_24050_7150# a_2475_7174# a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X629 VDD rowon_n[10] a_20946_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X630 a_25966_9158# row_n[7] a_26458_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X631 VDD rowon_n[4] a_32994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X632 a_26970_5142# row_n[3] a_27462_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X633 a_25966_18194# a_2275_18218# a_26058_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X634 a_30074_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X635 a_19942_8154# a_2275_8178# a_20034_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X636 VDD VSS a_30986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X637 VSS row_n[0] a_10298_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X638 a_31078_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X639 a_20946_4138# a_2275_4162# a_21038_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X640 VDD VDD a_19942_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X641 a_5278_14218# rowon_n[12] a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X642 a_15318_14218# rowon_n[12] a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X643 a_30074_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X644 a_20338_15222# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X645 a_2475_17214# a_1957_17214# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X646 a_12402_5504# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X647 a_13006_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X648 VSS row_n[2] a_4274_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X649 a_13310_17230# rowon_n[15] a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X650 a_6890_13174# a_2275_13198# a_6982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X651 a_16930_13174# a_2275_13198# a_17022_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X652 a_7286_7190# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X653 a_3270_17230# rowon_n[15] a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X654 a_29070_5142# a_2475_5166# a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X655 VSS row_n[11] a_4274_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X656 VSS row_n[11] a_14314_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X657 a_32082_12170# a_2475_12194# a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X658 a_11302_10202# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X659 a_19942_13174# row_n[11] a_20434_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X660 VSS row_n[4] a_21342_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X661 a_32994_12170# row_n[10] a_33486_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X662 a_14010_11166# a_2475_11190# a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X663 a_24962_6146# a_2275_6170# a_25054_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X664 a_31078_18194# a_2475_18218# a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X665 a_3970_11166# a_2475_11190# a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X666 a_2874_9158# a_2275_9182# a_2966_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X667 VDD rowon_n[5] a_17934_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X668 a_29982_7150# row_n[5] a_30474_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X669 a_35094_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X670 a_28978_2130# row_n[0] a_29470_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X671 a_31990_18194# VDD a_32482_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X672 VDD rowon_n[13] a_2874_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X673 VDD rowon_n[13] a_12914_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X674 vcm a_2275_14202# a_32082_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X675 a_10394_12532# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X676 a_4370_4500# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X677 a_14410_11528# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X678 a_18026_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X679 a_4370_11528# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X680 a_17022_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X681 VDD a_2161_5166# a_2275_5166# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X682 vcm a_2275_17214# a_30074_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X683 a_13918_5142# a_2275_5166# a_14010_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X684 a_33390_2170# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X685 a_14410_2492# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X686 VSS row_n[6] a_25358_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X687 VSS row_n[2] a_26362_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X688 a_35398_8194# rowon_n[6] a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X689 a_26058_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X690 a_35002_5142# row_n[3] a_35494_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X691 a_9994_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X692 VSS row_n[14] a_19334_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X693 a_23350_14218# rowon_n[12] a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X694 a_29374_12210# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X695 VSS row_n[9] a_20338_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X696 VSS row_n[8] a_33390_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X697 a_11302_4178# rowon_n[2] a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X698 a_24050_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X699 a_33998_11166# a_2275_11190# a_34090_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X700 a_10298_10202# rowon_n[8] a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X701 a_26458_4500# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X702 a_24962_13174# a_2275_13198# a_25054_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X703 a_17934_7150# a_2275_7174# a_18026_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X704 a_18938_3134# a_2275_3158# a_19030_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X705 VDD VDD a_17934_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X706 a_28466_14540# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X707 VDD rowon_n[10] a_31990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X708 a_28066_10162# a_2475_10186# a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X709 a_10998_5142# a_2475_5166# a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X710 a_20034_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X711 a_8990_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X712 VSS row_n[7] a_8290_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X713 a_28978_10162# row_n[8] a_29470_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X714 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X715 a_3270_3174# rowon_n[1] a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X716 VDD rowon_n[2] a_10906_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X717 VSS VDD a_34394_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X718 a_31382_15222# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X719 a_9902_10162# a_2275_10186# a_9994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X720 a_2161_8178# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X721 vcm a_2275_6170# a_23046_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X722 a_11302_18234# VDD a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X723 a_35398_14218# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X724 a_33086_6146# a_2475_6170# a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X725 a_29070_18194# a_2475_18218# a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X726 VSS row_n[12] a_12306_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X727 a_20338_5182# rowon_n[3] a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X728 a_30474_17552# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X729 vcm a_2275_15206# a_26058_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X730 a_30074_13174# a_2475_13198# a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X731 a_8386_9520# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X732 a_15014_7150# a_2475_7174# a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X733 a_25054_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X734 a_16018_3134# a_2475_3158# a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X735 a_24050_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X736 a_2874_17190# a_2275_17214# a_2966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X737 a_9994_17190# a_2475_17214# a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X738 a_12914_17190# a_2275_17214# a_13006_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X739 VDD VSS a_2874_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X740 a_34490_16548# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X741 a_30986_13174# row_n[11] a_31478_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X742 VDD rowon_n[6] a_21950_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X743 vcm a_2275_5166# a_12002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X744 VDD rowon_n[14] a_10906_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X745 vcm a_2275_10186# a_17022_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X746 a_9902_8154# row_n[6] a_10394_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X747 a_8290_1166# VSS a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X748 VSS row_n[2] a_34394_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X749 a_6890_14178# row_n[12] a_7382_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X750 a_16930_14178# row_n[12] a_17422_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X751 vcm a_2275_10186# a_6982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X752 a_8990_9158# a_2475_9182# a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X753 VDD rowon_n[1] a_19942_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X754 vcm a_2275_4162# a_28066_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X755 a_24354_7190# rowon_n[5] a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X756 a_2475_6170# a_1957_6170# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X757 a_7986_2130# a_2475_2154# a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X758 a_25358_3174# rowon_n[1] a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X759 a_29070_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X760 a_13310_3174# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X761 a_15318_9198# rowon_n[7] a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X762 a_32994_9158# a_2275_9182# a_33086_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X763 a_32082_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X764 VDD rowon_n[4] a_26970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X765 vcm a_2275_3158# a_17022_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X766 a_34490_4500# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X767 vcm a_2275_18218# a_7986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X768 vcm a_2275_18218# a_18026_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X769 VSS row_n[15] a_26362_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X770 a_30378_15222# rowon_n[13] a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X771 vcm a_2275_7174# a_16018_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X772 a_14922_6146# row_n[4] a_15414_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X773 a_31990_2130# a_2275_2154# a_32082_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X774 a_34394_14218# rowon_n[12] a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X775 a_27366_13214# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X776 VSS row_n[9] a_31382_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X777 VDD VSS a_24962_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X778 a_22042_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X779 a_12914_1126# VDD a_13406_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X780 VSS row_n[3] a_19334_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X781 a_13006_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X782 a_35094_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X783 a_5278_2170# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X784 a_29374_5182# rowon_n[3] a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X785 a_2966_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X786 a_22954_14178# a_2275_14202# a_23046_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X787 VDD rowon_n[7] a_14922_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X788 a_7286_8194# rowon_n[6] a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X789 a_18330_1166# en_bit_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15 M=2
X790 VDD VDD a_28978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X791 a_6982_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X792 a_17022_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X793 a_26458_15544# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X794 VDD rowon_n[11] a_29982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X795 a_26058_11166# a_2475_11190# a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X796 vcm a_2275_2154# a_8990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X797 a_30378_10202# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X798 VDD a_2161_12194# a_2275_12194# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X799 a_26970_11166# row_n[9] a_27462_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X800 a_23046_1126# a_2475_1150# a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X801 a_19430_3496# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X802 a_22042_5142# a_2475_5166# a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X803 VDD rowon_n[1] a_28978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X804 a_24962_14178# row_n[12] a_25454_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X805 vcm a_2275_10186# a_25054_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X806 a_23958_7150# row_n[5] a_24450_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X807 a_8990_12170# a_2475_12194# a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X808 a_28370_9198# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X809 a_19334_16226# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X810 vcm a_2275_16210# a_24050_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X811 a_21950_2130# row_n[0] a_22442_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X812 a_10906_18194# a_2275_18218# a_10998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X813 a_18026_18194# a_2475_18218# a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X814 a_9294_16226# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X815 a_7986_18194# a_2475_18218# a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X816 a_9390_12532# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X817 a_2475_11190# a_1957_11190# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X818 a_27366_2170# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X819 a_33390_3174# rowon_n[1] a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X820 a_10998_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X821 a_18426_18556# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X822 a_27062_3134# a_2475_3158# a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X823 a_8386_18556# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X824 vcm a_2275_9182# a_31078_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X825 a_17326_8194# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X826 a_3970_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X827 a_27974_9158# row_n[7] a_28466_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X828 a_28978_5142# row_n[3] a_29470_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X829 a_6890_8154# row_n[6] a_7382_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X830 VSS row_n[0] a_12306_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X831 a_22954_4138# a_2275_4162# a_23046_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X832 a_32082_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X833 VDD VSS a_32994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X834 a_33086_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X835 a_2161_17214# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X836 a_28370_15222# rowon_n[13] a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X837 VSS row_n[10] a_25358_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X838 a_30074_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X839 a_14410_5504# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X840 a_2966_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X841 VSS row_n[9] a_29374_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X842 a_15014_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X843 a_16018_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X844 a_9294_7190# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X845 VDD rowon_n[12] a_23958_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X846 a_12002_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X847 a_34090_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X848 a_10906_7150# a_2275_7174# a_10998_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X849 a_11910_3134# a_2275_3158# a_12002_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X850 a_9294_10202# rowon_n[8] a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X851 VSS row_n[4] a_23350_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X852 a_33086_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X853 VDD rowon_n[11] a_27974_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X854 a_25454_10524# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X855 a_10998_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X856 a_23350_17230# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X857 a_33998_14178# a_2275_14202# a_34090_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X858 a_4882_9158# a_2275_9182# a_4974_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X859 VDD rowon_n[0] a_17934_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X860 a_2161_18218# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X861 a_29982_2130# row_n[0] a_30474_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X862 a_3878_2130# a_2275_2154# a_3970_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X863 VSS row_n[13] a_7286_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X864 VSS row_n[13] a_17326_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X865 a_22042_15182# a_2475_15206# a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X866 a_4274_12210# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X867 a_14314_12210# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X868 a_15926_5142# a_2275_5166# a_16018_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X869 a_16930_1126# a_2275_1150# a_17022_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X870 a_18330_11206# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X871 vcm a_2275_11190# a_23046_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X872 a_35398_2170# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X873 VSS row_n[2] a_28370_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X874 a_22954_15182# row_n[13] a_23446_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X875 a_17022_13174# a_2475_13198# a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X876 a_8290_11206# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X877 VSS row_n[6] a_27366_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X878 a_6982_13174# a_2475_13198# a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X879 a_9902_13174# a_2275_13198# a_9994_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X880 a_1957_4162# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X881 VDD rowon_n[15] a_5886_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X882 VDD rowon_n[15] a_15926_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X883 a_3366_14540# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X884 a_13406_14540# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X885 a_17422_13536# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X886 a_13918_10162# row_n[8] a_14410_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X887 a_2161_2154# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X888 a_7382_13536# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X889 a_3878_10162# row_n[8] a_4370_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X890 vcm a_2275_8178# a_20034_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X891 vcm a_2275_4162# a_21038_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X892 a_13310_4178# rowon_n[2] a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X893 a_26970_9158# a_2275_9182# a_27062_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X894 a_30074_8154# a_2475_8178# a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X895 VSS row_n[5] a_16322_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X896 a_31078_4138# a_2475_4162# a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X897 a_28466_4500# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X898 a_6378_7512# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X899 a_13006_5142# a_2475_5166# a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X900 a_22042_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X901 a_22346_17230# rowon_n[15] a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X902 vcm a_2275_15206# a_10998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X903 VDD rowon_n[4] a_19942_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X904 a_4882_18194# VDD a_5374_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X905 a_14922_18194# VDD a_15414_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X906 a_26362_16226# rowon_n[14] a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X907 vcm a_2275_14202# a_4974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X908 vcm a_2275_14202# a_15014_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X909 VSS row_n[11] a_23350_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X910 a_8990_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X911 VDD rowon_n[2] a_12914_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X912 vcm a_2275_6170# a_25054_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X913 a_35094_6146# a_2475_6170# a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X914 a_27974_15182# a_2275_15206# a_28066_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X915 a_32082_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X916 vcm a_2275_9182# a_2966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X917 VDD rowon_n[13] a_21950_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X918 a_17326_11206# rowon_n[9] a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X919 a_11302_1166# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X920 a_22346_5182# rowon_n[3] a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X921 VDD rowon_n[12] a_35002_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X922 a_7286_11206# rowon_n[9] a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X923 a_17022_7150# a_2475_7174# a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X924 a_10298_5182# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X925 a_27062_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X926 a_18026_3134# a_2475_3158# a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X927 a_23446_11528# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X928 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X929 a_21342_18234# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X930 VDD rowon_n[6] a_23958_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X931 vcm a_2275_5166# a_14010_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X932 a_34394_17230# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X933 VDD rowon_n[1] a_21950_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X934 VSS row_n[15] a_11302_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X935 a_9902_3134# row_n[1] a_10394_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X936 a_29982_18194# a_2275_18218# a_30074_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X937 VSS row_n[14] a_15318_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X938 a_20034_16186# a_2475_16210# a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X939 a_12306_13214# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X940 vcm a_2275_17214# a_29070_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X941 VSS row_n[14] a_5278_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X942 a_10998_15182# a_2475_15206# a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X943 a_33086_15182# a_2475_15206# a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X944 a_21342_9198# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X945 VSS row_n[7] a_31382_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X946 a_26362_7190# rowon_n[5] a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X947 a_9994_2130# a_2475_2154# a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X948 a_27366_3174# rowon_n[1] a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X949 a_15318_3174# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X950 a_20946_16186# row_n[14] a_21438_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X951 a_5278_6186# rowon_n[4] a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X952 a_33998_15182# row_n[13] a_34490_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X953 a_15014_14178# a_2475_14202# a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X954 vcm a_2275_11190# a_34090_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X955 a_17326_9198# rowon_n[7] a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X956 a_35002_9158# a_2275_9182# a_35094_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X957 a_19430_6508# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X958 VDD VDD a_13918_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X959 a_11398_15544# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X960 a_4974_14178# a_2475_14202# a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X961 vcm a_2275_7174# a_18026_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X962 VDD rowon_n[4] a_28978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X963 vcm a_2275_3158# a_19030_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X964 VDD VDD a_3878_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X965 a_20034_3134# a_2475_3158# a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X966 a_11910_11166# row_n[9] a_12402_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X967 a_33998_2130# a_2275_2154# a_34090_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X968 VDD VSS a_26970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X969 a_20946_9158# row_n[7] a_21438_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X970 a_26058_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X971 a_14922_1126# VDD a_15414_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X972 a_21950_5142# row_n[3] a_22442_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X973 a_31478_9520# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X974 a_2475_14202# a_1957_14202# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X975 a_9902_14178# row_n[12] a_10394_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X976 vcm a_2275_10186# a_9994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X977 a_21342_12210# rowon_n[10] a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X978 VDD rowon_n[7] a_16930_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X979 a_9294_8194# rowon_n[6] a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X980 a_20338_18234# VDD a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X981 a_31382_1166# VSS a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X982 a_17022_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X983 a_25054_1126# a_2475_1150# a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X984 VSS row_n[12] a_21342_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X985 a_6982_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X986 a_24050_5142# a_2475_5166# a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X987 a_21950_17190# a_2275_17214# a_22042_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X988 VDD rowon_n[8] a_20946_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X989 a_25966_7150# row_n[5] a_26458_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X990 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X991 a_25966_16186# a_2275_16210# a_26058_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X992 a_30074_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X993 a_19942_6146# a_2275_6170# a_20034_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X994 a_9994_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X995 VDD rowon_n[14] a_19942_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X996 a_30074_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X997 a_23958_2130# row_n[0] a_24450_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X998 a_20338_13214# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X999 a_33390_12210# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1000 a_2475_15206# a_1957_15206# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X1001 a_12002_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1002 a_29374_2170# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1003 a_13006_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1004 a_3270_15222# rowon_n[13] a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1005 a_13310_15222# rowon_n[13] a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1006 VSS row_n[10] a_10298_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1007 a_7286_5182# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1008 a_32386_18234# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1009 a_19334_8194# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1010 a_29070_3134# a_2475_3158# a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1011 a_32482_14540# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1012 vcm a_2275_12194# a_28066_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1013 VSS row_n[9] a_4274_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1014 VSS row_n[9] a_14314_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1015 a_32082_10162# a_2475_10186# a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1016 vcm a_2275_9182# a_33086_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1017 a_19942_11166# row_n[9] a_20434_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1018 a_8898_8154# row_n[6] a_9390_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1019 VSS row_n[6] a_20338_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1020 VSS row_n[2] a_21342_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1021 vcm a_2275_18218# a_27062_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1022 a_31078_16186# a_2475_16210# a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1023 a_32994_10162# row_n[8] a_33486_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1024 a_30378_8194# rowon_n[6] a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1025 VSS row_n[0] a_14314_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1026 a_24962_4138# a_2275_4162# a_25054_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1027 a_34090_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1028 VDD rowon_n[3] a_17934_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1029 vcm a_2275_2154# a_32082_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1030 a_35094_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1031 a_29982_5142# row_n[3] a_30474_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1032 a_31990_16186# row_n[14] a_32482_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1033 VDD rowon_n[11] a_2874_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1034 VDD rowon_n[11] a_12914_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1035 a_10394_10524# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1036 a_4974_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1037 a_6890_3134# row_n[1] a_7382_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1038 a_17022_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1039 a_18026_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1040 a_2161_12194# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1041 VDD a_2161_3158# a_2275_3158# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X1042 a_13918_3134# a_2275_3158# a_14010_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1043 a_21438_4500# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1044 vcm a_2275_15206# a_30074_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1045 a_12914_7150# a_2275_7174# a_13006_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1046 VSS row_n[4] a_25358_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1047 VSS row_n[7] a_3270_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1048 a_35398_6186# rowon_n[4] a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1049 a_18330_18234# VDD a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1050 a_32386_12210# rowon_n[10] a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1051 VSS row_n[12] a_19334_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1052 a_29374_10202# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1053 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=2.7075 pd=21.85 as=0.2755 ps=2.19 w=1.9 l=0.22 M=2
X1054 a_24050_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1055 a_20946_12170# a_2275_12194# a_21038_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1056 a_5886_2130# a_2275_2154# a_5978_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1057 a_18938_1126# a_2275_1150# a_19030_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1058 a_17934_5142# a_2275_5166# a_18026_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1059 VDD rowon_n[14] a_17934_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1060 a_28466_12532# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1061 VDD rowon_n[8] a_31990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1062 a_3366_9520# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1063 VSS row_n[6] a_29374_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1064 a_20034_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1065 a_10998_3134# a_2475_3158# a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1066 a_8990_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1067 a_16418_8516# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1068 VSS row_n[15] a_30378_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1069 a_3270_1166# VSS a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1070 VSS row_n[14] a_34394_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1071 a_31382_13214# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1072 a_3970_9158# a_2475_9182# a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1073 a_32386_7190# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1074 a_2161_6170# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1075 a_11302_16226# rowon_n[14] a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1076 vcm a_2275_4162# a_23046_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1077 a_25054_17190# a_2475_17214# a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1078 a_28978_9158# a_2275_9182# a_29070_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1079 a_32082_8154# a_2475_8178# a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1080 VSS row_n[5] a_18330_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1081 a_33086_4138# a_2475_4162# a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1082 a_29070_16186# a_2475_16210# a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1083 vcm a_2275_13198# a_26058_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1084 a_2966_2130# a_2475_2154# a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1085 a_20338_3174# rowon_n[1] a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1086 VDD VDD a_32994_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1087 a_25966_17190# row_n[15] a_26458_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1088 a_30474_15544# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1089 a_30074_11166# a_2475_11190# a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1090 a_8386_7512# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1091 a_15014_5142# a_2475_5166# a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1092 a_16018_1126# a_2475_1150# a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1093 a_24050_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1094 a_2874_15182# a_2275_15206# a_2966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1095 a_9994_15182# a_2475_15206# a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1096 a_12914_15182# a_2275_15206# a_13006_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1097 a_10298_9198# rowon_n[7] a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1098 a_30986_11166# row_n[9] a_31478_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1099 VDD rowon_n[4] a_21950_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1100 a_6378_2492# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1101 vcm a_2275_3158# a_12002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1102 vcm a_2275_7174# a_10998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1103 a_9902_6146# row_n[4] a_10394_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1104 a_6890_12170# row_n[10] a_7382_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1105 a_16930_12170# row_n[10] a_17422_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1106 VDD en_bit_n[0] a_19942_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1107 vcm a_2275_9182# a_4974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1108 a_25358_1166# VSS a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1109 a_2475_4162# a_1957_4162# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X1110 a_24354_5182# rowon_n[3] a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1111 VDD rowon_n[7] a_9902_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1112 a_13310_1166# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1113 a_29070_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1114 vcm a_2275_17214# a_14010_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1115 a_27974_10162# a_2275_10186# a_28066_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1116 vcm a_2275_2154# a_3970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1117 vcm a_2275_17214# a_3970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1118 VDD rowon_n[6] a_25966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1119 vcm a_2275_1150# a_17022_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1120 a_29374_18234# VDD a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1121 vcm a_2275_16210# a_7986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1122 vcm a_2275_16210# a_18026_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1123 VSS row_n[13] a_26362_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1124 a_30378_13214# rowon_n[11] a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1125 vcm a_2275_5166# a_16018_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1126 a_27366_11206# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1127 VDD rowon_n[1] a_23958_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1128 a_22042_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1129 VSS row_n[1] a_19334_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1130 VDD rowon_n[15] a_24962_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1131 a_13006_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1132 a_35094_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1133 a_31990_12170# a_2275_12194# a_32082_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1134 a_23350_9198# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1135 a_28370_7190# rowon_n[5] a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1136 a_29374_3174# rowon_n[1] a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1137 a_2966_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1138 VSS row_n[7] a_33390_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1139 VDD rowon_n[5] a_14922_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1140 a_7286_6186# rowon_n[4] a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1141 VDD rowon_n[14] a_28978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1142 a_6982_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1143 a_17022_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1144 a_26458_13536# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1145 VDD rowon_n[9] a_29982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1146 vcm a_2275_9182# a_27062_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1147 a_22346_2170# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1148 VDD a_2161_10186# a_2275_10186# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X1149 a_24050_12170# a_2475_12194# a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1150 a_19430_1488# en_bit_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1151 a_22042_3134# a_2475_3158# a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1152 VSS row_n[10] a_9294_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1153 a_12306_8194# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1154 a_28066_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1155 VDD VSS a_28978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1156 VSS VDD a_18330_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1157 a_23046_18194# a_2475_18218# a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1158 a_24962_12170# row_n[10] a_25454_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1159 a_22954_9158# row_n[7] a_23446_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1160 a_23958_5142# row_n[3] a_24450_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1161 VSS VDD a_8290_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1162 a_8990_10162# a_2475_10186# a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1163 a_33486_9520# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1164 a_23958_18194# VDD a_24450_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1165 a_19334_14218# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1166 vcm a_2275_14202# a_24050_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1167 a_10906_16186# a_2275_16210# a_10998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1168 a_18026_16186# a_2475_16210# a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1169 VDD rowon_n[12] a_7894_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1170 a_9294_14218# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1171 a_7986_16186# a_2475_16210# a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1172 a_9390_10524# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1173 a_33390_1166# VSS a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1174 a_10998_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1175 a_18426_16548# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1176 a_4274_7190# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1177 a_27062_1126# a_2475_1150# a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1178 a_8386_16548# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1179 a_17326_6186# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1180 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1181 a_27974_7150# row_n[5] a_28466_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1182 vcm a_2275_12194# a_13006_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1183 a_6890_6146# row_n[4] a_7382_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1184 vcm a_2275_12194# a_2966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1185 a_32082_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1186 a_25966_2130# row_n[0] a_26458_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1187 a_2161_15206# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1188 a_28370_13214# rowon_n[11] a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1189 VSS row_n[8] a_25358_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1190 vcm a_2275_18218# a_12002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1191 a_25966_11166# a_2275_11190# a_26058_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1192 a_14010_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1193 a_15014_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1194 a_9294_5182# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1195 VDD rowon_n[10] a_23958_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1196 vcm a_2275_9182# a_35094_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1197 a_10906_5142# a_2275_5166# a_10998_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1198 a_11910_1126# a_2275_1150# a_12002_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1199 a_30378_2170# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1200 a_18330_2170# rowon_n[0] a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1201 VSS row_n[2] a_23350_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1202 a_28978_18194# a_2275_18218# a_29070_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1203 a_33086_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1204 VDD rowon_n[9] a_27974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1205 VSS row_n[6] a_22346_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1206 a_32386_8194# rowon_n[6] a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1207 a_10998_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1208 vcm a_2275_2154# a_34090_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1209 a_23350_15222# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1210 a_26058_8154# a_2475_8178# a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1211 a_8898_3134# row_n[1] a_9390_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1212 a_6982_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1213 a_16322_17230# rowon_n[15] a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1214 a_6282_17230# rowon_n[15] a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1215 a_2161_16210# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1216 a_21950_9158# a_2275_9182# a_22042_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1217 VSS row_n[5] a_11302_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1218 a_22442_17552# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1219 VSS row_n[11] a_7286_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1220 VSS row_n[11] a_17326_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1221 a_22042_13174# a_2475_13198# a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1222 a_35094_12170# a_2475_12194# a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1223 a_4274_10202# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1224 a_14314_10202# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1225 a_14922_7150# a_2275_7174# a_15014_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1226 a_15926_3134# a_2275_3158# a_16018_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1227 a_23446_4500# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1228 a_2966_12170# a_2475_12194# a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1229 a_13006_12170# a_2475_12194# a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1230 a_22954_13174# row_n[11] a_23446_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1231 a_17022_11166# a_2475_11190# a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1232 VSS row_n[4] a_27366_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1233 a_6982_11166# a_2475_11190# a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1234 VSS row_n[7] a_5278_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1235 a_1957_18218# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1236 VDD rowon_n[13] a_5886_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1237 VDD rowon_n[13] a_15926_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1238 a_3366_12532# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1239 a_13406_12532# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1240 a_17422_11528# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1241 a_7382_11528# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1242 vcm a_2275_6170# a_20034_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1243 a_15318_18234# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1244 vcm a_2275_18218# a_20034_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1245 a_30074_6146# a_2475_6170# a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1246 VSS row_n[3] a_16322_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1247 a_7894_2130# a_2275_2154# a_7986_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1248 a_5278_18234# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1249 vcm a_2275_17214# a_33086_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1250 a_5374_9520# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1251 a_31990_8154# row_n[6] a_32482_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1252 a_6378_5504# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1253 a_24050_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1254 a_18426_8516# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1255 a_12002_7150# a_2475_7174# a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1256 a_22042_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1257 a_13006_3134# a_2475_3158# a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1258 a_10906_17190# row_n[15] a_11398_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1259 a_22346_15222# rowon_n[13] a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1260 vcm a_2275_13198# a_10998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1261 a_4882_16186# row_n[14] a_5374_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1262 a_14922_16186# row_n[14] a_15414_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1263 a_26362_14218# rowon_n[12] a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1264 VSS row_n[9] a_23350_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1265 a_16418_3496# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1266 a_34394_7190# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1267 vcm a_2275_4162# a_25054_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1268 a_27062_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1269 a_34090_8154# a_2475_8178# a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1270 a_35094_4138# a_2475_4162# a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1271 a_27974_13174# a_2275_13198# a_28066_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1272 a_1957_9182# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1273 VDD rowon_n[11] a_21950_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1274 a_21342_7190# rowon_n[5] a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1275 a_4974_2130# a_2475_2154# a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1276 a_22346_3174# rowon_n[1] a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1277 a_10298_3174# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1278 VDD rowon_n[10] a_35002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1279 a_17022_5142# a_2475_5166# a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1280 a_18026_1126# a_2475_1150# a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1281 a_12306_9198# rowon_n[7] a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1282 a_29982_9158# a_2275_9182# a_30074_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1283 a_21342_16226# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1284 vcm a_2275_7174# a_13006_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1285 VDD rowon_n[4] a_23958_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1286 a_8386_2492# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1287 vcm a_2275_3158# a_14010_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1288 a_34394_15222# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1289 a_12914_10162# a_2275_10186# a_13006_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1290 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1291 a_2874_10162# a_2275_10186# a_2966_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1292 VDD VSS a_21950_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1293 a_4274_18234# VDD a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1294 a_14314_18234# VDD a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1295 VSS row_n[13] a_11302_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1296 a_21038_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1297 a_9902_1126# VDD a_10394_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1298 a_20434_18556# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1299 a_29982_16186# a_2275_16210# a_30074_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1300 VSS row_n[12] a_15318_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1301 a_20034_14178# a_2475_14202# a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1302 a_12306_11206# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1303 a_33486_17552# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1304 vcm a_2275_15206# a_29070_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1305 VSS row_n[12] a_5278_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1306 a_10998_13174# a_2475_13198# a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1307 a_33086_13174# a_2475_13198# a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1308 a_15318_1166# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1309 a_27366_1166# VSS a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1310 a_26362_5182# rowon_n[3] a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1311 a_5886_17190# a_2275_17214# a_5978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1312 a_15926_17190# a_2275_17214# a_16018_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1313 VDD rowon_n[7] a_11910_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1314 a_4274_8194# rowon_n[6] a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1315 a_5278_4178# rowon_n[2] a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1316 VDD rowon_n[15] a_9902_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1317 a_33998_13174# row_n[11] a_34490_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1318 vcm a_2275_2154# a_5978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1319 VDD rowon_n[14] a_13918_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1320 a_11398_13536# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1321 VDD rowon_n[6] a_27974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1322 vcm a_2275_5166# a_18026_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1323 vcm a_2275_1150# a_19030_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1324 VDD rowon_n[14] a_3878_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1325 a_20034_1126# a_2475_1150# a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1326 a_20946_7150# row_n[5] a_21438_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1327 a_26058_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1328 VDD rowon_n[1] a_25966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1329 vcm a_2275_18218# a_31078_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1330 a_31478_7512# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1331 VDD rowon_n[2] a_4882_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1332 a_9902_12170# row_n[10] a_10394_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1333 a_21342_10202# rowon_n[8] a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1334 a_25358_9198# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1335 a_22042_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1336 VSS row_n[7] a_35398_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1337 VDD rowon_n[5] a_16930_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1338 a_9294_6186# rowon_n[4] a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1339 a_13006_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1340 a_35094_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1341 vcm a_2275_9182# a_29070_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1342 a_20338_16226# rowon_n[14] a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1343 a_2966_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1344 a_24354_2170# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1345 VDD rowon_n[0] a_14922_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1346 a_14314_8194# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1347 a_24050_3134# a_2475_3158# a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1348 a_25054_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1349 a_21950_15182# a_2275_15206# a_22042_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1350 a_24962_9158# row_n[7] a_25454_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1351 a_25966_5142# row_n[3] a_26458_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1352 a_16018_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1353 a_35494_9520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1354 a_3878_8154# row_n[6] a_4370_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1355 a_5978_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1356 a_25966_14178# a_2275_14202# a_26058_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1357 a_19942_4138# a_2275_4162# a_20034_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1358 a_9994_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1359 a_30074_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1360 a_20338_11206# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1361 a_33390_10202# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1362 a_2475_13198# a_1957_13198# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X1363 a_12002_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1364 a_13006_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1365 a_3270_13214# rowon_n[11] a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1366 a_13310_13214# rowon_n[11] a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1367 VSS row_n[8] a_10298_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1368 a_6282_7190# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1369 a_7286_3174# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1370 a_32386_16226# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1371 a_10906_11166# a_2275_11190# a_10998_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1372 a_19334_6186# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1373 a_29070_1126# a_2475_1150# a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1374 a_27974_14178# row_n[12] a_28466_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1375 a_32482_12532# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1376 vcm a_2275_10186# a_28066_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1377 a_14922_12170# a_2275_12194# a_15014_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1378 a_8898_6146# row_n[4] a_9390_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1379 VSS row_n[4] a_20338_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1380 vcm a_2275_16210# a_27062_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1381 a_31078_14178# a_2475_14202# a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1382 a_4882_12170# a_2275_12194# a_4974_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1383 a_30378_6186# rowon_n[4] a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1384 a_13918_18194# a_2275_18218# a_14010_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1385 a_31478_18556# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1386 a_34090_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1387 a_27974_2130# row_n[0] a_28466_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1388 a_3878_18194# a_2275_18218# a_3970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1389 VDD rowon_n[9] a_2874_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1390 VDD rowon_n[9] a_12914_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1391 a_6890_1126# VDD a_7382_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1392 a_17022_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1393 a_2161_10186# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1394 VDD a_2161_1150# a_2275_1150# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X1395 a_13918_1126# a_2275_1150# a_14010_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1396 a_29982_17190# row_n[15] a_30474_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1397 vcm a_2275_13198# a_30074_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1398 a_12914_5142# a_2275_5166# a_13006_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1399 VSS row_n[6] a_24354_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1400 VSS row_n[2] a_25358_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1401 a_11398_8516# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1402 a_34394_8194# rowon_n[6] a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1403 a_35398_4178# rowon_n[2] a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1404 a_18330_16226# rowon_n[14] a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1405 VSS row_n[10] a_28370_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1406 a_33086_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1407 a_32386_10202# rowon_n[8] a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1408 a_28066_8154# a_2475_8178# a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1409 a_8990_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1410 a_10998_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1411 a_24050_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1412 a_19030_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1413 VDD rowon_n[12] a_26970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1414 a_15014_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1415 a_23958_9158# a_2275_9182# a_24050_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1416 VSS row_n[5] a_13310_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1417 a_4974_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1418 a_17934_3134# a_2275_3158# a_18026_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1419 VDD rowon_n[2] a_35002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1420 a_25454_4500# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1421 a_28466_10524# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1422 a_3366_7512# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1423 VSS row_n[4] a_29374_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1424 a_10998_1126# a_2475_1150# a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1425 VSS row_n[7] a_7286_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1426 a_16418_6508# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1427 a_33390_18234# VDD a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1428 a_26362_17230# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1429 VSS row_n[13] a_30378_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1430 VSS row_n[12] a_34394_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1431 a_31382_11206# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1432 VSS row_n[0] a_6282_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1433 a_2161_4162# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1434 a_32386_5182# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1435 a_35002_17190# a_2275_17214# a_35094_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1436 a_11302_14218# rowon_n[12] a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1437 a_1957_13198# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1438 a_25054_15182# a_2475_15206# a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1439 a_7286_12210# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1440 a_17326_12210# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1441 vcm a_2275_12194# a_22042_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1442 a_32082_6146# a_2475_6170# a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1443 VSS row_n[3] a_18330_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1444 a_29070_14178# a_2475_14202# a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1445 vcm a_2275_11190# a_26058_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1446 a_33998_8154# row_n[6] a_34490_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1447 a_20338_1166# en_bit_n[0] a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1448 a_29470_18556# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1449 VDD rowon_n[14] a_32994_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1450 a_25966_15182# row_n[13] a_26458_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1451 a_30474_13536# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1452 a_7382_9520# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1453 a_8386_5504# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1454 a_24050_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1455 a_15014_3134# a_2475_3158# a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1456 a_2874_13174# a_2275_13198# a_2966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1457 a_9994_13174# a_2475_13198# a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1458 a_12914_13174# a_2275_13198# a_13006_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1459 a_14010_7150# a_2475_7174# a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1460 VDD rowon_n[15] a_8898_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1461 a_6378_14540# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1462 a_16418_14540# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1463 VDD rowon_n[6] a_20946_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1464 vcm a_2275_1150# a_12002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1465 a_31990_3134# row_n[1] a_32482_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1466 vcm a_2275_5166# a_10998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1467 a_18426_3496# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1468 a_6890_10162# row_n[8] a_7382_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1469 a_16930_10162# row_n[8] a_17422_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1470 a_23350_7190# rowon_n[5] a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1471 a_6982_2130# a_2475_2154# a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1472 a_24354_3174# rowon_n[1] a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1473 VDD rowon_n[5] a_9902_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1474 a_25358_17230# rowon_n[15] a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1475 vcm a_2275_15206# a_14010_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1476 vcm a_2275_15206# a_3970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1477 a_14314_9198# rowon_n[7] a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1478 vcm a_2275_9182# a_22042_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1479 VDD rowon_n[4] a_25966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1480 a_17934_18194# VDD a_18426_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1481 a_29374_16226# rowon_n[14] a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1482 vcm a_2275_14202# a_7986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1483 vcm a_2275_14202# a_18026_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1484 VSS row_n[11] a_26362_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1485 a_30378_11206# rowon_n[9] a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1486 vcm a_2275_7174# a_15014_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1487 vcm a_2275_3158# a_16018_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1488 a_7894_18194# VDD a_8386_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1489 a_30986_2130# a_2275_2154# a_31078_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1490 a_23046_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1491 VDD VSS a_23958_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1492 a_22042_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1493 VDD rowon_n[13] a_24962_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1494 a_13006_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1495 a_35094_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1496 a_29374_1166# VSS a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1497 a_28370_5182# rowon_n[3] a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1498 a_2966_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1499 a_25358_12210# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1500 VDD rowon_n[7] a_13918_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1501 VDD rowon_n[3] a_14922_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1502 a_7286_4178# rowon_n[2] a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1503 a_26458_11528# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1504 a_29982_11166# a_2275_11190# a_30074_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1505 a_6282_8194# rowon_n[6] a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1506 vcm a_2275_2154# a_7986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1507 a_24354_18234# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1508 a_24450_14540# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1509 a_24050_10162# a_2475_10186# a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1510 a_2475_9182# a_1957_9182# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X1511 a_22042_1126# a_2475_1150# a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1512 VSS row_n[8] a_9294_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1513 a_12306_6186# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1514 a_28066_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1515 VDD rowon_n[1] a_27974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1516 a_32994_18194# a_2275_18218# a_33086_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1517 VSS row_n[14] a_18330_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1518 a_23046_16186# a_2475_16210# a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1519 a_24962_10162# row_n[8] a_25454_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1520 a_22954_7150# row_n[5] a_23446_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1521 VSS row_n[14] a_8290_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1522 a_33486_7512# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1523 VDD rowon_n[2] a_6890_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1524 a_23958_16186# row_n[14] a_24450_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1525 a_20946_2130# row_n[0] a_21438_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1526 a_10906_14178# a_2275_14202# a_10998_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1527 a_18026_14178# a_2475_14202# a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1528 VDD rowon_n[10] a_7894_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1529 a_31478_2492# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1530 VDD VDD a_16930_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1531 a_7986_14178# a_2475_14202# a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1532 VDD VDD a_6890_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1533 a_26362_2170# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1534 VDD rowon_n[0] a_16930_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1535 a_4274_5182# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1536 vcm a_2275_9182# a_30074_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1537 a_16322_8194# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1538 a_17326_4178# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1539 a_27974_5142# row_n[3] a_28466_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1540 vcm a_2275_10186# a_13006_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1541 a_5886_8154# row_n[6] a_6378_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1542 a_2874_14178# row_n[12] a_3366_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1543 a_12914_14178# row_n[12] a_13406_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1544 a_24354_12210# rowon_n[10] a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1545 vcm a_2275_10186# a_2966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1546 a_21950_10162# a_2275_10186# a_22042_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1547 a_32082_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1548 a_28370_11206# rowon_n[9] a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1549 a_21038_8154# a_2475_8178# a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1550 a_3878_3134# row_n[1] a_4370_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1551 vcm a_2275_16210# a_12002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1552 a_14010_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1553 a_15014_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1554 a_16930_4138# row_n[2] a_17422_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1555 a_9994_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1556 a_8290_7190# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1557 a_9294_3174# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1558 VDD rowon_n[8] a_23958_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1559 a_9902_7150# a_2275_7174# a_9994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1560 a_10906_3134# a_2275_3158# a_10998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1561 VSS row_n[15] a_22346_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1562 a_28978_16186# a_2275_16210# a_29070_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1563 a_33086_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1564 VSS row_n[4] a_22346_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1565 a_32386_6186# rowon_n[4] a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1566 a_10998_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1567 a_23350_13214# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1568 a_26058_6146# a_2475_6170# a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1569 a_8898_1126# VDD a_9390_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1570 a_16322_15222# rowon_n[13] a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1571 VSS row_n[10] a_13310_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1572 a_6282_15222# rowon_n[13] a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1573 a_2161_14202# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1574 VSS row_n[10] a_3270_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1575 VSS row_n[3] a_11302_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1576 a_2874_2130# a_2275_2154# a_2966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1577 a_22442_15544# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1578 a_35494_14540# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1579 VSS row_n[9] a_7286_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1580 VSS row_n[9] a_17326_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1581 a_22042_11166# a_2475_11190# a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1582 a_35094_10162# a_2475_10186# a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1583 a_14922_5142# a_2275_5166# a_15014_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1584 a_15926_1126# a_2275_1150# a_16018_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1585 a_22954_11166# row_n[9] a_23446_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1586 a_2966_10162# a_2475_10186# a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1587 a_13006_10162# a_2475_10186# a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1588 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1589 VSS row_n[2] a_27366_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1590 VDD rowon_n[12] a_11910_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1591 a_13406_8516# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1592 VDD rowon_n[11] a_5886_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1593 VDD rowon_n[11] a_15926_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1594 a_3366_10524# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1595 a_13406_10524# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1596 a_11302_17230# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1597 a_11398_3496# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1598 vcm a_2275_4162# a_20034_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1599 a_15318_16226# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1600 vcm a_2275_16210# a_20034_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1601 a_25966_9158# a_2275_9182# a_26058_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1602 VSS row_n[5] a_15318_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1603 VSS row_n[1] a_16322_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1604 a_30074_4138# a_2475_4162# a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1605 a_14010_18194# a_2475_18218# a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1606 a_5278_16226# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1607 vcm a_2275_15206# a_33086_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1608 a_27462_4500# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1609 a_3970_18194# a_2475_18218# a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1610 a_5374_7512# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1611 a_31990_6146# row_n[4] a_32482_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1612 a_5978_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1613 a_18426_6508# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1614 a_12002_5142# a_2475_5166# a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1615 a_13006_1126# a_2475_1150# a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1616 a_14410_18556# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1617 a_10906_15182# row_n[13] a_11398_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1618 a_22346_13214# rowon_n[11] a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1619 vcm a_2275_11190# a_10998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1620 VSS row_n[7] a_9294_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1621 a_4370_18556# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1622 a_35398_12210# rowon_n[10] a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1623 a_3366_2492# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1624 a_16418_1488# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1625 a_27062_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1626 a_23958_12170# a_2275_12194# a_24050_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1627 VSS row_n[0] a_8290_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1628 a_34394_5182# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1629 a_34090_6146# a_2475_6170# a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1630 a_1957_7174# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1631 VDD rowon_n[9] a_21950_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1632 a_9390_9520# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1633 a_10298_1166# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1634 a_22346_1166# VSS a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1635 a_21342_5182# rowon_n[3] a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1636 VDD rowon_n[8] a_35002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1637 a_17022_3134# a_2475_3158# a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1638 VSS VDD a_20338_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1639 VSS row_n[15] a_33390_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1640 a_33998_3134# row_n[1] a_34490_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1641 a_21342_14218# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1642 VDD rowon_n[6] a_22954_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1643 a_6890_7150# a_2275_7174# a_6982_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1644 vcm a_2275_5166# a_13006_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1645 vcm a_2275_1150# a_14010_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1646 a_10298_17230# rowon_n[15] a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1647 a_34394_13214# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1648 a_28066_17190# a_2475_17214# a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1649 a_4274_16226# rowon_n[14] a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1650 a_14314_16226# rowon_n[14] a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1651 VSS row_n[11] a_11302_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1652 a_21038_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1653 VDD rowon_n[1] a_20946_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1654 a_20434_16548# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1655 a_29982_14178# a_2275_14202# a_30074_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1656 a_28978_17190# row_n[15] a_29470_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1657 a_33486_15544# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1658 vcm a_2275_13198# a_29070_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1659 a_10998_11166# a_2475_11190# a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1660 a_33086_11166# a_2475_11190# a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1661 a_20338_9198# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1662 a_8990_2130# a_2475_2154# a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1663 a_26362_3174# rowon_n[1] a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1664 a_5886_15182# a_2275_15206# a_5978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1665 a_15926_15182# a_2275_15206# a_16018_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1666 VSS row_n[7] a_30378_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1667 VDD rowon_n[5] a_11910_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1668 a_4274_6186# rowon_n[4] a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1669 VDD rowon_n[13] a_9902_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1670 a_33998_11166# row_n[9] a_34490_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1671 a_16322_9198# rowon_n[7] a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1672 vcm a_2275_9182# a_24050_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1673 a_19030_7150# a_2475_7174# a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1674 a_10298_12210# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1675 a_11398_11528# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1676 VDD rowon_n[4] a_27974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1677 VDD rowon_n[0] a_9902_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1678 vcm a_2275_3158# a_18026_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1679 VDD VSS a_25966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1680 a_32994_2130# a_2275_2154# a_33086_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1681 a_15318_2170# rowon_n[0] a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1682 a_26058_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1683 a_19942_9158# row_n[7] a_20434_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1684 a_25054_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1685 a_20946_5142# row_n[3] a_21438_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1686 vcm a_2275_16210# a_31078_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1687 a_30474_9520# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1688 a_31478_5504# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1689 a_9902_10162# row_n[8] a_10394_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1690 vcm a_2275_17214# a_17022_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1691 VDD rowon_n[7] a_15926_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1692 a_8290_8194# rowon_n[6] a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1693 VDD rowon_n[3] a_16930_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1694 a_9294_4178# rowon_n[2] a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1695 vcm a_2275_17214# a_6982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1696 a_20338_14218# rowon_n[12] a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1697 a_21038_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1698 a_14314_6186# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1699 a_24050_1126# a_2475_1150# a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1700 a_25054_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1701 a_21950_13174# a_2275_13198# a_22042_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1702 a_24962_7150# row_n[5] a_25454_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1703 a_16018_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1704 a_35494_7512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1705 a_3878_6146# row_n[4] a_4370_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1706 a_5978_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1707 VDD rowon_n[2] a_8898_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1708 a_9994_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1709 VSS row_n[10] a_32386_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1710 a_22954_2130# row_n[0] a_23446_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1711 a_33486_2492# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1712 VSS VDD a_31382_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1713 a_2475_11190# a_1957_11190# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X1714 a_28370_2170# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1715 a_12002_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1716 VDD rowon_n[12] a_30986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1717 a_27062_12170# a_2475_12194# a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1718 a_3270_11206# rowon_n[9] a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1719 a_13310_11206# rowon_n[9] a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1720 a_6282_5182# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1721 a_7286_1166# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1722 a_32386_14218# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1723 a_19334_4178# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1724 a_26058_18194# a_2475_18218# a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1725 a_27974_12170# row_n[10] a_28466_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1726 a_32482_10524# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1727 a_18330_8194# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1728 VSS row_n[2] a_20338_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1729 a_26970_18194# VDD a_27462_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1730 a_30378_17230# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1731 vcm a_2275_14202# a_27062_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1732 a_7894_8154# row_n[6] a_8386_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1733 a_30378_4178# rowon_n[2] a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1734 a_13918_16186# a_2275_16210# a_14010_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1735 a_31478_16548# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1736 vcm a_2275_2154# a_31078_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1737 a_34090_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1738 a_3878_16186# a_2275_16210# a_3970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1739 a_23046_8154# a_2475_8178# a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1740 a_3970_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1741 a_5886_3134# row_n[1] a_6378_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1742 a_17022_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1743 vcm a_2275_17214# a_25054_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1744 a_18938_4138# row_n[2] a_19430_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1745 vcm a_2275_11190# a_30074_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1746 a_20434_4500# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1747 a_29982_15182# row_n[13] a_30474_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1748 a_12914_3134# a_2275_3158# a_13006_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1749 VDD rowon_n[2] a_29982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1750 vcm a_2275_12194# a_16018_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1751 VSS row_n[4] a_24354_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1752 vcm a_2275_12194# a_5978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1753 a_11398_6508# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1754 a_34394_6186# rowon_n[4] a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1755 a_18330_14218# rowon_n[12] a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1756 VSS row_n[8] a_28370_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1757 a_19030_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1758 a_28978_11166# a_2275_11190# a_29070_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1759 a_28066_6146# a_2475_6170# a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1760 a_20034_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1761 a_19030_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1762 VDD rowon_n[10] a_26970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1763 VSS row_n[3] a_13310_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1764 a_4882_2130# a_2275_2154# a_4974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1765 a_17934_1126# a_2275_1150# a_18026_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1766 a_3366_5504# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1767 VSS row_n[2] a_29374_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1768 a_15414_8516# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1769 a_16018_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1770 VSS VDD a_29374_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1771 a_33390_16226# rowon_n[14] a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1772 a_26362_15222# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1773 VSS row_n[11] a_30378_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1774 VSS a_2161_6170# a_2275_6170# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X1775 a_13406_3496# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1776 a_19334_7190# rowon_n[5] a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1777 a_31382_7190# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1778 a_32386_3174# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1779 a_9294_17230# rowon_n[15] a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1780 a_35002_15182# a_2275_15206# a_35094_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1781 a_25454_17552# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1782 a_21950_14178# row_n[12] a_22442_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1783 a_25054_13174# a_2475_13198# a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1784 a_7286_10202# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1785 a_17326_10202# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1786 vcm a_2275_10186# a_22042_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1787 a_27974_9158# a_2275_9182# a_28066_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1788 VSS row_n[5] a_17326_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1789 VSS row_n[1] a_18330_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1790 a_32082_4138# a_2475_4162# a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1791 a_5978_12170# a_2475_12194# a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1792 a_16018_12170# a_2475_12194# a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1793 a_33998_6146# row_n[4] a_34490_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1794 a_29470_4500# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1795 a_29470_16548# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1796 a_25966_13174# row_n[11] a_26458_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1797 a_30474_11528# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1798 a_7382_7512# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1799 a_7986_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1800 a_14010_5142# a_2475_5166# a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1801 a_15014_1126# a_2475_1150# a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1802 a_9994_11166# a_2475_11190# a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1803 a_26970_2130# a_2275_2154# a_27062_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1804 VDD rowon_n[13] a_8898_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1805 a_6378_12532# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1806 a_16418_12532# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1807 VDD rowon_n[4] a_20946_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1808 a_31990_1126# VDD a_32482_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1809 a_5374_2492# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1810 vcm a_2275_3158# a_10998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1811 vcm a_2275_7174# a_9994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1812 a_18426_1488# en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1813 a_16930_8154# a_2275_8178# a_17022_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1814 a_18330_18234# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1815 vcm a_2275_18218# a_23046_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1816 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1817 a_8290_18234# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1818 a_24354_1166# VSS a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1819 a_23350_5182# rowon_n[3] a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1820 a_27062_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1821 VDD rowon_n[3] a_9902_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1822 a_13918_17190# row_n[15] a_14410_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1823 a_25358_15222# rowon_n[13] a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1824 vcm a_2275_13198# a_14010_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1825 a_2161_9182# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1826 vcm a_2275_2154# a_2966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1827 a_3878_17190# row_n[15] a_4370_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1828 vcm a_2275_13198# a_3970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1829 vcm a_2275_1150# a_16018_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1830 a_17934_16186# row_n[14] a_18426_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1831 a_29374_14218# rowon_n[12] a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1832 VSS row_n[9] a_26362_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1833 a_8898_7150# a_2275_7174# a_8990_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1834 vcm a_2275_5166# a_15014_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1835 a_7894_16186# row_n[14] a_8386_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1836 a_31078_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1837 a_23046_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1838 VDD rowon_n[1] a_22954_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1839 VDD rowon_n[11] a_24962_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1840 a_28370_3174# rowon_n[1] a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1841 a_25358_10202# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1842 VSS row_n[7] a_32386_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1843 VDD rowon_n[5] a_13918_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1844 a_6282_6186# rowon_n[4] a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1845 a_24354_16226# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1846 vcm a_2275_9182# a_26058_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1847 a_8290_12210# rowon_n[10] a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1848 a_15926_10162# a_2275_10186# a_16018_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1849 VSS row_n[0] a_31382_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1850 a_21342_2170# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1851 VDD rowon_n[0] a_11910_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1852 a_24450_12532# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1853 a_5886_10162# a_2275_10186# a_5978_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1854 a_2475_7174# a_1957_7174# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X1855 a_5978_7150# a_2475_7174# a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1856 a_7286_18234# VDD a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1857 a_17326_18234# VDD a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1858 a_11302_8194# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1859 a_27062_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1860 a_35002_2130# a_2275_2154# a_35094_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1861 VDD VSS a_27974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1862 a_17326_2170# rowon_n[0] a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1863 a_28066_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1864 a_12306_4178# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1865 a_23446_18556# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1866 a_32994_16186# a_2275_16210# a_33086_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1867 VSS row_n[12] a_18330_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1868 a_23046_14178# a_2475_14202# a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1869 a_22954_5142# row_n[3] a_23446_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1870 VSS row_n[12] a_8290_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1871 a_32482_9520# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1872 a_33486_5504# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1873 a_18938_17190# a_2275_17214# a_19030_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1874 a_8898_17190# a_2275_17214# a_8990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1875 VDD rowon_n[8] a_7894_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1876 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1877 VDD rowon_n[14] a_16930_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1878 VDD rowon_n[14] a_6890_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1879 a_11910_4138# row_n[2] a_12402_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1880 vcm a_2275_12194# a_35094_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1881 a_3270_7190# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1882 a_4274_3174# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1883 a_16322_6186# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1884 vcm a_2275_18218# a_34090_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1885 vcm a_2275_7174# a_6982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1886 a_12914_12170# row_n[10] a_13406_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1887 a_5886_6146# row_n[4] a_6378_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1888 a_2874_12170# row_n[10] a_3366_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1889 a_25054_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1890 a_24354_10202# rowon_n[8] a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1891 a_16018_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1892 a_21038_6146# a_2475_6170# a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1893 a_35494_2492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1894 a_3878_1126# en_C0_n a_4370_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1895 a_24962_2130# row_n[0] a_25454_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1896 a_11910_18194# VDD a_12402_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1897 vcm a_2275_14202# a_12002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1898 a_5978_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1899 VDD rowon_n[12] a_18938_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1900 a_29070_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1901 a_14010_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1902 a_8290_5182# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1903 a_9294_1166# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1904 a_28066_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1905 vcm a_2275_17214# a_9994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1906 a_9902_5142# a_2275_5166# a_9994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1907 a_10906_1126# a_2275_1150# a_10998_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1908 VSS row_n[2] a_22346_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1909 VSS row_n[13] a_22346_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1910 a_28978_14178# a_2275_14202# a_29070_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1911 a_32386_4178# rowon_n[2] a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1912 a_31382_8194# rowon_n[6] a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1913 vcm a_2275_2154# a_33086_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1914 a_23350_11206# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1915 a_25054_8154# a_2475_8178# a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1916 a_26058_4138# a_2475_4162# a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1917 a_7894_3134# row_n[1] a_8386_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1918 VDD rowon_n[15] a_20946_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1919 a_16322_13214# rowon_n[11] a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1920 VSS row_n[8] a_13310_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1921 a_6282_13214# rowon_n[11] a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1922 a_3878_11166# a_2275_11190# a_3970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1923 a_13918_11166# a_2275_11190# a_14010_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1924 VSS row_n[8] a_3270_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1925 a_20946_9158# a_2275_9182# a_21038_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1926 VSS row_n[5] a_10298_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1927 VSS row_n[1] a_11302_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1928 a_22442_13536# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1929 a_35494_12532# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1930 a_31078_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1931 a_14922_3134# a_2275_3158# a_15014_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1932 a_22442_4500# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1933 a_17934_12170# a_2275_12194# a_18026_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1934 VDD rowon_n[2] a_31990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1935 a_7894_12170# a_2275_12194# a_7986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1936 VDD rowon_n[10] a_11910_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1937 a_13406_6508# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1938 VSS row_n[7] a_4274_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1939 a_6890_18194# a_2275_18218# a_6982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1940 a_16930_18194# a_2275_18218# a_17022_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1941 VDD rowon_n[9] a_5886_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1942 VDD rowon_n[9] a_15926_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1943 VSS VDD a_14314_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1944 a_11302_15222# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1945 a_11398_1488# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1946 VSS VDD a_4274_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1947 a_32082_17190# a_2475_17214# a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1948 VSS row_n[0] a_3270_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1949 a_19942_18194# VDD a_20434_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1950 a_15318_14218# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1951 vcm a_2275_14202# a_20034_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1952 VSS row_n[3] a_15318_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1953 VSS VDD a_16322_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1954 a_32994_17190# row_n[15] a_33486_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1955 a_14010_16186# a_2475_16210# a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1956 a_5278_14218# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1957 vcm a_2275_13198# a_33086_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1958 a_10394_17552# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1959 a_3970_16186# a_2475_16210# a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1960 a_4370_9520# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1961 VDD rowon_n[6] a_18938_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1962 a_30986_8154# row_n[6] a_31478_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1963 a_5374_5504# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1964 a_17422_8516# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1965 a_5978_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1966 a_12002_3134# a_2475_3158# a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1967 a_14410_16548# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1968 a_10906_13174# row_n[11] a_11398_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1969 a_22346_11206# rowon_n[9] a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1970 a_18026_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1971 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0.2755 pd=2.19 as=0.551 ps=4.38 w=1.9 l=0.22 M=4
X1972 a_4370_16548# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1973 a_35398_10202# rowon_n[8] a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1974 a_15414_3496# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1975 a_27062_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1976 VSS row_n[7] a_26362_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1977 a_33390_7190# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1978 a_34394_3174# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1979 a_18026_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1980 a_34090_4138# a_2475_4162# a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1981 a_7986_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1982 a_1957_5166# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1983 a_9390_7512# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1984 a_3970_2130# a_2475_2154# a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1985 a_21342_3174# rowon_n[1] a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1986 a_35002_10162# a_2275_10186# a_35094_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1987 a_9994_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1988 a_17022_1126# a_2475_1150# a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1989 a_29374_17230# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1990 VSS row_n[14] a_20338_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1991 VSS row_n[13] a_33390_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1992 a_11302_9198# rowon_n[7] a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1993 a_28978_2130# a_2275_2154# a_29070_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1994 VDD rowon_n[4] a_22954_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1995 a_6890_5142# a_2275_5166# a_6982_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1996 a_7382_2492# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1997 vcm a_2275_3158# a_13006_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1998 a_10298_15222# rowon_n[13] a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1999 a_34394_11206# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2000 a_26458_9520# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2001 a_18938_8154# a_2275_8178# a_19030_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2002 a_24962_18194# a_2275_18218# a_25054_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2003 VDD VSS a_20946_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2004 a_10298_2170# rowon_n[0] a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2005 a_21038_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2006 VDD rowon_n[15] a_31990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2007 a_28066_15182# a_2475_15206# a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2008 a_4274_14218# rowon_n[12] a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2009 a_14314_14218# rowon_n[12] a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2010 VSS row_n[9] a_11302_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2011 a_20034_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2012 a_28978_15182# row_n[13] a_29470_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2013 a_33486_13536# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2014 vcm a_2275_11190# a_29070_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2015 VDD rowon_n[3] a_11910_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2016 a_26362_1166# VSS a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2017 a_5886_13174# a_2275_13198# a_5978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2018 a_15926_13174# a_2275_13198# a_16018_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2019 VDD rowon_n[7] a_10906_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2020 a_3270_8194# rowon_n[6] a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2021 a_4274_4178# rowon_n[2] a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2022 VDD rowon_n[11] a_9902_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2023 vcm a_2275_2154# a_4974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2024 a_19030_5142# a_2475_5166# a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2025 a_10298_10202# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2026 vcm a_2275_1150# a_18026_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2027 a_30074_18194# a_2475_18218# a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2028 a_16018_8154# a_2475_8178# a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2029 a_19942_7150# row_n[5] a_20434_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2030 a_25054_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2031 a_30986_18194# VDD a_31478_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2032 vcm a_2275_14202# a_31078_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2033 a_30474_7512# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2034 VDD rowon_n[2] a_3878_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2035 vcm a_2275_15206# a_17022_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2036 VSS row_n[7] a_34394_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2037 VDD rowon_n[5] a_15926_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2038 a_8290_6186# rowon_n[4] a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2039 vcm a_2275_15206# a_6982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2040 vcm a_2275_9182# a_28066_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2041 a_23350_2170# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2042 VDD rowon_n[0] a_13918_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2043 a_21038_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2044 VSS row_n[0] a_33390_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2045 a_25358_8194# rowon_n[6] a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2046 a_7986_7150# a_2475_7174# a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2047 a_14314_4178# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2048 VSS a_2161_16210# a_2275_16210# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X2049 a_25054_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2050 a_13310_8194# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2051 a_29070_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2052 vcm a_2275_2154# a_27062_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2053 a_24962_5142# row_n[3] a_25454_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2054 a_16018_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2055 a_34490_9520# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2056 a_35494_5504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2057 a_5978_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2058 a_28370_12210# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2059 VSS row_n[8] a_32386_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2060 a_2874_8154# row_n[6] a_3366_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2061 vcm a_2275_8178# a_17022_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2062 a_32994_11166# a_2275_11190# a_33086_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2063 a_31990_7150# a_2275_7174# a_32082_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2064 a_27366_18234# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2065 VSS row_n[14] a_31382_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2066 a_12002_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2067 a_27462_14540# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2068 VDD rowon_n[10] a_30986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2069 a_27062_10162# a_2475_10186# a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2070 a_6282_3174# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2071 a_13918_4138# row_n[2] a_14410_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2072 a_5278_7190# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2073 a_26058_16186# a_2475_16210# a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2074 a_27974_10162# row_n[8] a_28466_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2075 a_18330_6186# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2076 VDD VDD a_29982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2077 vcm a_2275_7174# a_8990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2078 a_26970_16186# row_n[14] a_27462_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2079 a_30378_15222# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2080 a_7894_6146# row_n[4] a_8386_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2081 VDD a_2161_17214# a_2275_17214# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X2082 a_13918_14178# a_2275_14202# a_14010_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2083 a_3878_14178# a_2275_14202# a_3970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2084 a_23046_6146# a_2475_6170# a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2085 a_5886_1126# VDD a_6378_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2086 vcm a_2275_15206# a_25054_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2087 a_8990_17190# a_2475_17214# a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2088 a_29982_13174# row_n[11] a_30474_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2089 a_12914_1126# a_2275_1150# a_13006_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2090 vcm a_2275_10186# a_16018_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2091 VSS row_n[2] a_24354_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2092 a_9390_17552# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2093 a_5886_14178# row_n[12] a_6378_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2094 a_15926_14178# row_n[12] a_16418_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2095 a_27366_12210# rowon_n[10] a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2096 vcm a_2275_10186# a_5978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2097 a_10394_8516# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2098 a_10998_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2099 a_33390_8194# rowon_n[6] a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2100 a_27366_7190# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2101 a_34394_4178# rowon_n[2] a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2102 vcm a_2275_2154# a_35094_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2103 a_19030_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2104 a_27062_8154# a_2475_8178# a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2105 a_28066_4138# a_2475_4162# a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2106 a_19030_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2107 VDD rowon_n[8] a_26970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2108 a_22954_9158# a_2275_9182# a_23046_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2109 VSS row_n[5] a_12306_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2110 VSS row_n[1] a_13310_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2111 a_33086_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2112 VDD rowon_n[2] a_33998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2113 a_24450_4500# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2114 VSS row_n[15] a_25358_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2115 a_2966_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2116 a_15414_6508# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2117 a_16018_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2118 a_21950_2130# a_2275_2154# a_22042_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2119 VSS row_n[14] a_29374_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2120 a_33390_14218# rowon_n[12] a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2121 a_26362_13214# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2122 VSS row_n[9] a_30378_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2123 VSS a_2161_4162# a_2275_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X2124 a_13406_1488# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2125 a_12002_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2126 a_34090_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2127 VSS row_n[10] a_16322_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2128 a_21038_12170# a_2475_12194# a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2129 a_11910_8154# a_2275_8178# a_12002_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2130 a_32386_1166# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2131 a_31382_5182# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2132 a_19334_5182# rowon_n[3] a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2133 a_9294_15222# rowon_n[13] a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2134 a_35002_13174# a_2275_13198# a_35094_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2135 VSS row_n[10] a_6282_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2136 VSS row_n[0] a_5278_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2137 VDD VDD a_27974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2138 a_25454_15544# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2139 a_21950_12170# row_n[10] a_22442_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2140 a_25054_11166# a_2475_11190# a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2141 VSS row_n[3] a_17326_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2142 a_5978_10162# a_2475_10186# a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2143 a_16018_10162# a_2475_10186# a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2144 VDD rowon_n[12] a_14922_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2145 a_25966_11166# row_n[9] a_26458_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2146 a_32994_8154# row_n[6] a_33486_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2147 a_7382_5504# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2148 a_7986_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2149 a_14010_3134# a_2475_3158# a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2150 VDD rowon_n[12] a_4882_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2151 VDD rowon_n[11] a_8898_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2152 a_6378_10524# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2153 a_16418_10524# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2154 vcm a_2275_1150# a_10998_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2155 a_30986_3134# row_n[1] a_31478_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2156 VDD rowon_n[1] a_18938_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2157 a_14314_17230# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2158 a_3878_7150# a_2275_7174# a_3970_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2159 vcm a_2275_5166# a_9994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2160 a_4274_17230# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2161 a_16930_6146# a_2275_6170# a_17022_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2162 a_17422_3496# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2163 a_18330_16226# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2164 vcm a_2275_16210# a_23046_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2165 VSS row_n[7] a_28370_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2166 a_35398_7190# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2167 a_9902_18194# a_2275_18218# a_9994_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2168 a_17022_18194# a_2475_18218# a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2169 a_8290_16226# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2170 a_1957_9182# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2171 a_6982_18194# a_2475_18218# a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2172 a_23350_3174# rowon_n[1] a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2173 a_17422_18556# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2174 a_13918_15182# row_n[13] a_14410_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2175 a_25358_13214# rowon_n[11] a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2176 a_1957_12194# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2177 vcm a_2275_11190# a_14010_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2178 a_2161_7174# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2179 a_7382_18556# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2180 a_3878_15182# row_n[13] a_4370_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2181 vcm a_2275_11190# a_3970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2182 a_13310_9198# rowon_n[7] a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2183 vcm a_2275_9182# a_21038_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2184 a_31078_9158# a_2475_9182# a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2185 a_8898_5142# a_2275_5166# a_8990_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2186 a_9390_2492# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2187 vcm a_2275_3158# a_15014_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2188 a_28466_9520# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2189 a_26970_12170# a_2275_12194# a_27062_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2190 a_22042_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2191 VDD VSS a_22954_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2192 a_29982_2130# a_2275_2154# a_30074_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2193 a_12306_2170# rowon_n[0] a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2194 a_23046_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2195 VSS row_n[10] a_24354_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2196 VDD rowon_n[9] a_24962_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2197 a_28370_1166# VSS a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2198 VDD rowon_n[7] a_12914_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2199 VDD rowon_n[3] a_13918_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2200 a_6282_4178# rowon_n[2] a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2201 VSS VDD a_23350_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2202 VDD rowon_n[12] a_22954_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2203 a_24354_14218# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2204 a_19030_12170# a_2475_12194# a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2205 a_8290_10202# rowon_n[8] a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2206 a_32082_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2207 a_24450_10524# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2208 a_2475_5166# a_1957_5166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X2209 a_5978_5142# a_2475_5166# a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2210 a_7286_16226# rowon_n[14] a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2211 a_17326_16226# rowon_n[14] a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2212 a_18026_8154# a_2475_8178# a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2213 a_11302_6186# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2214 a_27062_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2215 a_23446_16548# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2216 a_32994_14178# a_2275_14202# a_33086_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2217 a_32482_7512# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2218 VDD rowon_n[2] a_5886_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2219 a_18938_15182# a_2275_15206# a_19030_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2220 a_8898_15182# a_2275_15206# a_8990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2221 a_30474_2492# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2222 a_19942_2130# row_n[0] a_20434_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2223 a_3270_12210# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2224 a_13310_12210# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2225 a_25358_2170# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2226 VDD rowon_n[0] a_15926_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2227 a_12306_18234# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2228 a_35002_14178# row_n[12] a_35494_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2229 vcm a_2275_10186# a_35094_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2230 a_27366_8194# rowon_n[6] a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2231 a_9994_7150# a_2475_7174# a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2232 a_3270_5182# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2233 VSS row_n[0] a_35398_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2234 a_4274_1166# en_C0_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15 M=2
X2235 a_15318_8194# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2236 vcm a_2275_2154# a_29070_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2237 a_16322_4178# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2238 vcm a_2275_16210# a_34090_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2239 a_12402_14540# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2240 a_21038_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2241 vcm a_2275_5166# a_6982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2242 a_12914_10162# row_n[8] a_13406_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2243 a_4882_8154# row_n[6] a_5374_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2244 VSS a_2161_11190# a_2275_11190# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X2245 a_2874_10162# row_n[8] a_3366_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2246 vcm a_2275_8178# a_19030_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2247 a_20034_8154# a_2475_8178# a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2248 a_21038_4138# a_2475_4162# a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2249 a_11910_16186# row_n[14] a_12402_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2250 a_33998_7150# a_2275_7174# a_34090_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2251 a_2874_3134# row_n[1] a_3366_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2252 VDD rowon_n[10] a_18938_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2253 a_14010_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2254 a_8290_3174# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2255 a_15926_4138# row_n[2] a_16418_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2256 a_21342_17230# rowon_n[15] a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2257 a_28066_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2258 vcm a_2275_15206# a_9994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2259 a_9902_3134# a_2275_3158# a_9994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2260 VSS row_n[11] a_22346_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2261 a_31382_6186# rowon_n[4] a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2262 VSS row_n[10] a_35398_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2263 a_12306_12210# rowon_n[10] a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2264 a_25054_6146# a_2475_6170# a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2265 a_7894_1126# VDD a_8386_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2266 VDD rowon_n[13] a_20946_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2267 a_6282_11206# rowon_n[9] a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2268 a_16322_11206# rowon_n[9] a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2269 a_26970_8154# row_n[6] a_27462_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2270 VDD rowon_n[12] a_33998_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2271 VSS row_n[3] a_10298_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2272 VSS VDD a_11302_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2273 a_22442_11528# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2274 a_35494_10524# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2275 a_14922_1126# a_2275_1150# a_15014_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2276 a_20338_18234# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2277 a_33390_17230# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2278 VDD rowon_n[8] a_11910_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2279 a_12402_8516# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2280 a_13006_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2281 a_29374_7190# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2282 VSS row_n[15] a_10298_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2283 a_6890_16186# a_2275_16210# a_6982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2284 a_16930_16186# a_2275_16210# a_17022_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2285 a_29070_8154# a_2475_8178# a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2286 VSS row_n[14] a_14314_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2287 a_11302_13214# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2288 a_10394_3496# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2289 vcm a_2275_17214# a_28066_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2290 VSS row_n[14] a_4274_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2291 a_32082_15182# a_2475_15206# a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2292 VSS row_n[7] a_21342_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2293 a_19942_16186# row_n[14] a_20434_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2294 a_19030_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2295 VSS row_n[1] a_15318_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2296 a_32994_15182# row_n[13] a_33486_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2297 a_14010_14178# a_2475_14202# a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2298 vcm a_2275_11190# a_33086_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2299 a_24962_9158# a_2275_9182# a_25054_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2300 a_35094_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2301 VSS row_n[5] a_14314_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2302 vcm a_2275_7174# a_32082_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2303 VDD VDD a_12914_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2304 a_10394_15544# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2305 a_3970_14178# a_2475_14202# a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2306 a_4370_7512# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2307 VDD rowon_n[4] a_18938_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2308 a_30986_6146# row_n[4] a_31478_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2309 VDD VDD a_2874_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2310 vcm a_2275_12194# a_8990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2311 vcm a_2275_12194# a_19030_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2312 a_4974_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2313 a_17422_6508# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2314 a_12002_1126# a_2475_1150# a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2315 a_5978_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2316 a_10906_11166# row_n[9] a_11398_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2317 VDD a_2161_8178# a_2275_8178# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X2318 a_18026_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2319 a_23958_2130# a_2275_2154# a_24050_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2320 a_23046_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2321 a_21438_9520# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2322 a_13918_8154# a_2275_8178# a_14010_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2323 a_15414_1488# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2324 VSS row_n[0] a_7286_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2325 a_33390_5182# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2326 a_1957_3158# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2327 a_32386_17230# rowon_n[15] a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2328 a_35002_8154# row_n[6] a_35494_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2329 a_9390_5504# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2330 a_21342_1166# VSS a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2331 a_9994_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2332 a_29374_15222# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2333 VSS row_n[12] a_20338_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2334 VSS row_n[11] a_33390_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2335 a_20946_17190# a_2275_17214# a_21038_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2336 a_5886_7150# a_2275_7174# a_5978_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2337 vcm a_2275_1150# a_13006_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2338 a_32994_3134# row_n[1] a_33486_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2339 a_6890_3134# a_2275_3158# a_6982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2340 a_10298_13214# rowon_n[11] a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2341 a_26458_7512# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2342 a_18938_6146# a_2275_6170# a_19030_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2343 a_24962_16186# a_2275_16210# a_25054_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2344 a_8990_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2345 a_28466_17552# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2346 VDD rowon_n[13] a_31990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2347 a_28066_13174# a_2475_13198# a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2348 a_10998_8154# a_2475_8178# a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2349 a_20034_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2350 a_11910_12170# a_2275_12194# a_12002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2351 a_28978_13174# row_n[11] a_29470_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2352 a_33486_11528# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2353 VDD rowon_n[9] a_9902_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2354 VDD rowon_n[5] a_10906_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2355 a_3270_6186# rowon_n[4] a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2356 a_31382_18234# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2357 vcm a_2275_9182# a_23046_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2358 a_19030_3134# a_2475_3158# a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2359 a_33086_9158# a_2475_9182# a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2360 vcm a_2275_18218# a_26058_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2361 a_30074_16186# a_2475_16210# a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2362 a_20338_8194# rowon_n[6] a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2363 a_2966_7150# a_2475_7174# a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2364 a_24050_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2365 a_16018_6146# a_2475_6170# a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2366 vcm a_2275_2154# a_22042_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2367 a_14314_2170# rowon_n[0] a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2368 a_25054_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2369 a_19942_5142# row_n[3] a_20434_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2370 a_30986_16186# row_n[14] a_31478_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2371 a_30474_5504# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2372 vcm a_2275_8178# a_12002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2373 a_16930_17190# row_n[15] a_17422_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2374 vcm a_2275_13198# a_17022_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2375 VDD rowon_n[3] a_15926_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2376 a_8290_4178# rowon_n[2] a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2377 a_6890_17190# row_n[15] a_7382_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2378 vcm a_2275_13198# a_6982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2379 a_21038_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2380 a_2475_9182# a_1957_9182# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X2381 a_25358_6186# rowon_n[4] a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2382 a_7986_5142# a_2475_5166# a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2383 VSS a_2161_14202# a_2275_14202# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X2384 a_13310_6186# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2385 a_29070_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2386 a_31382_12210# rowon_n[10] a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2387 vcm a_2275_7174# a_3970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2388 a_34490_7512# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2389 a_2874_6146# row_n[4] a_3366_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2390 a_28370_10202# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2391 vcm a_2275_6170# a_17022_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2392 VDD rowon_n[2] a_7894_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2393 a_30378_18234# VDD a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2394 a_19942_12170# a_2275_12194# a_20034_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2395 a_32482_2492# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2396 a_31990_5142# a_2275_5166# a_32082_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2397 a_27366_16226# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2398 VSS row_n[12] a_31382_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2399 a_18938_10162# a_2275_10186# a_19030_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2400 a_31990_17190# a_2275_17214# a_32082_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2401 a_27462_12532# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2402 a_8898_10162# a_2275_10186# a_8990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2403 VDD rowon_n[8] a_30986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2404 VSS row_n[6] a_19334_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2405 a_6282_1166# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2406 a_29374_8194# rowon_n[6] a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2407 a_5278_5182# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2408 a_26058_14178# a_2475_14202# a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2409 a_18330_4178# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2410 a_26458_18556# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2411 VDD rowon_n[14] a_29982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2412 vcm a_2275_5166# a_8990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2413 a_30378_13214# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2414 a_22346_7190# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2415 VDD a_2161_15206# a_2275_15206# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X2416 vcm a_2275_2154# a_30074_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2417 VSS row_n[15] a_9294_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2418 a_24050_17190# a_2475_17214# a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2419 a_22042_8154# a_2475_8178# a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2420 a_4882_3134# row_n[1] a_5374_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2421 a_23046_4138# a_2475_4162# a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2422 vcm a_2275_13198# a_25054_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2423 a_24962_17190# row_n[15] a_25454_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2424 a_17934_4138# row_n[2] a_18426_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2425 a_8990_15182# a_2475_15206# a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2426 a_29982_11166# row_n[9] a_30474_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2427 a_9390_15544# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2428 a_5886_12170# row_n[10] a_6378_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2429 a_15926_12170# row_n[10] a_16418_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2430 a_28066_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2431 a_27366_10202# rowon_n[8] a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2432 a_10394_6508# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2433 a_10998_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2434 a_33390_6186# rowon_n[4] a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2435 a_27366_5182# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2436 a_19030_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2437 a_27062_6146# a_2475_6170# a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2438 a_28978_8154# row_n[6] a_29470_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2439 a_19030_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2440 vcm a_2275_17214# a_13006_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2441 VSS row_n[3] a_12306_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2442 VSS VDD a_13310_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2443 vcm a_2275_17214# a_2966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2444 a_26970_3134# row_n[1] a_27462_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2445 a_28370_18234# VDD a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2446 VSS row_n[13] a_25358_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2447 a_22346_12210# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2448 a_2966_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2449 a_14410_8516# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2450 a_16018_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2451 VSS row_n[12] a_29374_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2452 a_26362_11206# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2453 a_15014_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2454 VSS a_2161_2154# a_2275_2154# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X2455 VDD rowon_n[15] a_23958_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2456 a_12002_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2457 a_34090_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2458 a_21438_14540# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2459 a_30986_12170# a_2275_12194# a_31078_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2460 VSS row_n[8] a_16322_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2461 a_21038_10162# a_2475_10186# a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2462 a_18330_7190# rowon_n[5] a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2463 a_11910_6146# a_2275_6170# a_12002_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2464 a_31382_3174# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2465 a_19334_3174# rowon_n[1] a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2466 a_12402_3496# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2467 a_9294_13214# rowon_n[11] a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2468 a_6890_11166# a_2275_11190# a_6982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2469 a_16930_11166# a_2275_11190# a_17022_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2470 VSS row_n[8] a_6282_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2471 VSS row_n[7] a_23350_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2472 a_30378_7190# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2473 VDD rowon_n[14] a_27974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2474 a_25454_13536# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2475 a_21950_10162# row_n[8] a_22442_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2476 VSS row_n[1] a_17326_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2477 vcm a_2275_7174# a_34090_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2478 a_32994_6146# row_n[4] a_33486_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2479 VDD rowon_n[10] a_14922_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2480 a_14010_1126# a_2475_1150# a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2481 a_7986_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2482 VDD rowon_n[10] a_4882_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2483 a_6982_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2484 a_25966_2130# a_2275_2154# a_26058_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2485 VDD rowon_n[9] a_8898_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2486 VDD en_bit_n[2] a_18938_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2487 a_30986_1126# VDD a_31478_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2488 VSS VDD a_17326_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2489 a_22042_18194# a_2475_18218# a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2490 a_14314_15222# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2491 a_3878_5142# a_2275_5166# a_3970_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2492 a_4370_2492# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2493 vcm a_2275_3158# a_9994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2494 VSS VDD a_7286_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2495 a_13006_17190# a_2475_17214# a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2496 a_35094_17190# a_2475_17214# a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2497 a_4274_15222# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2498 a_23446_9520# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2499 a_15926_8154# a_2275_8178# a_16018_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2500 a_17422_1488# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2501 a_16930_4138# a_2275_4162# a_17022_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2502 a_22954_18194# VDD a_23446_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2503 a_2966_17190# a_2475_17214# a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2504 a_18330_14218# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2505 vcm a_2275_14202# a_23046_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2506 VSS row_n[0] a_9294_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2507 a_35398_5182# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2508 a_9902_16186# a_2275_16210# a_9994_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2509 a_17022_16186# a_2475_16210# a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2510 a_8290_14218# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2511 a_13406_17552# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2512 a_6982_16186# a_2475_16210# a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2513 a_23350_1166# VSS a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2514 a_3366_17552# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2515 a_17422_16548# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2516 a_13918_13174# row_n[11] a_14410_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2517 a_25358_11206# rowon_n[9] a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2518 a_1957_10186# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2519 a_2161_5166# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2520 a_7382_16548# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2521 a_3878_13174# row_n[11] a_4370_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2522 a_35002_3134# row_n[1] a_35494_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2523 a_7894_7150# a_2275_7174# a_7986_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2524 vcm a_2275_1150# a_15014_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2525 a_8898_3134# a_2275_3158# a_8990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2526 a_28466_7512# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2527 a_13006_8154# a_2475_8178# a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2528 a_22042_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2529 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0.551 pd=4.38 as=0.2755 ps=2.19 w=1.9 l=0.22 M=4
X2530 VSS row_n[8] a_24354_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2531 a_26458_2492# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2532 vcm a_2275_18218# a_10998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2533 a_24962_11166# a_2275_11190# a_25054_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2534 VDD rowon_n[5] a_12914_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2535 VSS row_n[14] a_23350_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2536 a_19430_14540# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2537 VDD rowon_n[10] a_22954_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2538 a_19030_10162# a_2475_10186# a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2539 vcm a_2275_9182# a_25054_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2540 a_35094_9158# a_2475_9182# a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2541 a_20338_2170# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2542 VDD rowon_n[0] a_10906_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2543 a_27974_18194# a_2275_18218# a_28066_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2544 a_32082_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2545 a_22346_8194# rowon_n[6] a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2546 a_4974_7150# a_2475_7174# a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2547 VSS row_n[0] a_30378_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2548 a_5978_3134# a_2475_3158# a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2549 a_2475_3158# a_1957_3158# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X2550 VDD VDD a_21950_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2551 VDD rowon_n[15] a_35002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2552 a_7286_14218# rowon_n[12] a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2553 a_17326_14218# rowon_n[12] a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2554 a_10298_8194# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2555 a_18026_6146# a_2475_6170# a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2556 vcm a_2275_2154# a_24050_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2557 a_16322_2170# rowon_n[0] a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2558 a_27062_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2559 a_11302_4178# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2560 a_32482_5504# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2561 a_8898_13174# a_2275_13198# a_8990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2562 a_18938_13174# a_2275_13198# a_19030_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2563 vcm a_2275_8178# a_14010_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2564 a_34090_12170# a_2475_12194# a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2565 a_3270_10202# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2566 a_13310_10202# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2567 a_12002_12170# a_2475_12194# a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2568 a_12306_16226# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2569 a_35002_12170# row_n[10] a_35494_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2570 a_27366_6186# rowon_n[4] a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2571 a_9994_5142# a_2475_5166# a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2572 a_3270_3174# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2573 a_10906_4138# row_n[2] a_11398_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2574 a_10998_18194# a_2475_18218# a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2575 a_33086_18194# a_2475_18218# a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2576 a_5278_9198# rowon_n[7] a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2577 a_15318_6186# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2578 a_33998_18194# VDD a_34490_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2579 vcm a_2275_14202# a_34090_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2580 a_12402_12532# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2581 a_19334_12210# rowon_n[10] a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2582 vcm a_2275_3158# a_6982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2583 vcm a_2275_7174# a_5978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2584 a_4882_6146# row_n[4] a_5374_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2585 a_11398_18556# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2586 vcm a_2275_6170# a_19030_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2587 a_20034_6146# a_2475_6170# a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2588 a_34490_2492# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2589 a_2874_1126# VDD a_3366_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2590 a_33998_5142# a_2275_5166# a_34090_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2591 VDD rowon_n[8] a_18938_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2592 a_21950_8154# row_n[6] a_22442_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2593 a_2475_17214# a_1957_17214# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X2594 VDD rowon_n[7] a_4882_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2595 a_8290_1166# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2596 a_9902_17190# row_n[15] a_10394_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2597 a_21342_15222# rowon_n[13] a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2598 a_28066_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2599 vcm a_2275_13198# a_9994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2600 a_9902_1126# a_2275_1150# a_9994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2601 VSS row_n[9] a_22346_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2602 a_31382_4178# rowon_n[2] a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2603 VSS row_n[8] a_35398_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2604 a_24354_7190# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2605 a_12306_10202# rowon_n[8] a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2606 a_24050_8154# a_2475_8178# a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2607 a_25054_4138# a_2475_4162# a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2608 VDD rowon_n[11] a_20946_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2609 a_26970_6146# row_n[4] a_27462_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2610 VDD rowon_n[10] a_33998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2611 VSS row_n[1] a_10298_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2612 a_19942_9158# a_2275_9182# a_20034_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2613 a_30074_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2614 a_20338_16226# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2615 VDD rowon_n[2] a_30986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2616 a_2475_18218# a_1957_18218# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X2617 a_33390_15222# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2618 a_12402_6508# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2619 a_16930_14178# a_2275_14202# a_17022_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2620 a_13006_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2621 a_29374_5182# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2622 a_3270_18234# VDD a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2623 a_13310_18234# VDD a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2624 VSS row_n[13] a_10298_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2625 a_6890_14178# a_2275_14202# a_6982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2626 a_7286_8194# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2627 a_29070_6146# a_2475_6170# a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2628 VSS row_n[12] a_14314_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2629 a_11302_11206# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2630 a_10394_1488# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2631 a_32482_17552# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2632 vcm a_2275_15206# a_28066_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2633 VSS row_n[12] a_4274_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2634 a_32082_13174# a_2475_13198# a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2635 a_4882_17190# a_2275_17214# a_4974_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2636 a_14922_17190# a_2275_17214# a_15014_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2637 VSS row_n[3] a_14314_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2638 VSS VDD a_15318_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2639 a_32994_13174# row_n[11] a_33486_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2640 a_28978_3134# row_n[1] a_29470_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2641 vcm a_2275_5166# a_32082_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2642 VDD rowon_n[14] a_12914_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2643 a_10394_13536# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2644 vcm a_2275_10186# a_19030_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2645 VDD rowon_n[6] a_17934_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2646 a_29982_8154# row_n[6] a_30474_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2647 a_4370_5504# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2648 VDD rowon_n[14] a_2874_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2649 a_8898_14178# row_n[12] a_9390_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2650 a_18938_14178# row_n[12] a_19430_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2651 vcm a_2275_10186# a_8990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2652 a_4974_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2653 a_5978_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2654 a_17022_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2655 VDD a_2161_6170# a_2275_6170# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X2656 a_18026_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2657 vcm a_2275_18218# a_30074_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2658 a_21438_7512# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2659 a_13918_6146# a_2275_6170# a_14010_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2660 a_14410_3496# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2661 a_33390_3174# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2662 VSS row_n[7] a_25358_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2663 a_35398_9198# rowon_n[7] a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2664 a_12002_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2665 a_34090_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2666 VSS row_n[15] a_28370_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2667 a_32386_15222# rowon_n[13] a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2668 a_35002_6146# row_n[4] a_35494_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2669 a_8990_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2670 a_9994_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2671 a_29374_13214# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2672 VSS row_n[9] a_33390_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2673 a_27974_2130# a_2275_2154# a_28066_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2674 a_24050_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2675 a_20946_15182# a_2275_15206# a_21038_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2676 a_5886_5142# a_2275_5166# a_5978_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2677 a_6890_1126# a_2275_1150# a_6982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2678 a_32994_1126# VDD a_33486_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2679 a_15014_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2680 a_10298_11206# rowon_n[9] a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2681 a_25454_9520# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2682 a_17934_8154# a_2275_8178# a_18026_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2683 a_18938_4138# a_2275_4162# a_19030_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2684 a_26458_5504# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2685 a_4974_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2686 a_24962_14178# a_2275_14202# a_25054_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2687 VDD rowon_n[7] a_35002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2688 a_8990_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2689 a_28466_15544# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2690 VDD rowon_n[11] a_31990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2691 a_28066_11166# a_2475_11190# a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2692 a_10998_6146# a_2475_6170# a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2693 a_20034_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2694 a_28978_11166# row_n[9] a_29470_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2695 a_9902_11166# a_2275_11190# a_9994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2696 a_2161_9182# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2697 VDD rowon_n[3] a_10906_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2698 a_3270_4178# rowon_n[2] a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2699 a_31382_16226# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2700 VSS row_n[5] a_6282_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2701 a_19030_1126# a_2475_1150# a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2702 vcm a_2275_17214# a_22042_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2703 a_7286_17230# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2704 a_17326_17230# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2705 vcm a_2275_16210# a_26058_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2706 a_30074_14178# a_2475_14202# a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2707 a_20338_6186# rowon_n[4] a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2708 a_2966_5142# a_2475_5166# a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2709 a_12914_18194# a_2275_18218# a_13006_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2710 a_30474_18556# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2711 a_15014_8154# a_2475_8178# a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2712 a_24050_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2713 a_16018_4138# a_2475_4162# a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2714 a_2874_18194# a_2275_18218# a_2966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2715 a_9994_18194# a_2475_18218# a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2716 a_28466_2492# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2717 vcm a_2275_6170# a_12002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2718 VDD rowon_n[2] a_2874_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2719 a_16930_15182# row_n[13] a_17422_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2720 vcm a_2275_11190# a_17022_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2721 a_6890_15182# row_n[13] a_7382_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2722 vcm a_2275_11190# a_6982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2723 VDD rowon_n[0] a_12914_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2724 VSS row_n[0] a_32386_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2725 a_24354_8194# rowon_n[6] a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2726 a_6982_7150# a_2475_7174# a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2727 a_7986_3134# a_2475_3158# a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2728 a_25358_4178# rowon_n[2] a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2729 VSS row_n[10] a_27366_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2730 vcm a_2275_2154# a_26058_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2731 a_29070_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2732 a_13310_4178# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2733 a_32082_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2734 a_31382_10202# rowon_n[8] a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2735 vcm a_2275_5166# a_3970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2736 a_34490_5504# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2737 vcm a_2275_8178# a_16018_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2738 vcm a_2275_4162# a_17022_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2739 VSS VDD a_26362_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2740 a_30378_16226# rowon_n[14] a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2741 VDD rowon_n[12] a_25966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2742 a_14010_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2743 a_30986_7150# a_2275_7174# a_31078_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2744 a_31990_3134# a_2275_3158# a_32082_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2745 a_27366_14218# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2746 a_3970_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2747 VDD rowon_n[2] a_24962_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2748 a_35094_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2749 a_31990_15182# a_2275_15206# a_32082_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2750 a_27462_10524# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2751 VSS row_n[4] a_19334_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2752 a_12914_4138# row_n[2] a_13406_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2753 a_2966_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2754 a_13006_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2755 a_29374_6186# rowon_n[4] a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2756 a_5278_3174# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2757 a_25358_17230# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2758 a_26458_16548# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2759 a_7286_9198# rowon_n[7] a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2760 vcm a_2275_7174# a_7986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2761 vcm a_2275_3158# a_8990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2762 a_30378_11206# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2763 a_22346_5182# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2764 VDD a_2161_13198# a_2275_13198# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X2765 VSS row_n[13] a_9294_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2766 a_24050_15182# a_2475_15206# a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2767 a_6282_12210# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2768 a_16322_12210# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2769 vcm a_2275_12194# a_21038_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2770 a_22042_6146# a_2475_6170# a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2771 a_4882_1126# VDD a_5374_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2772 vcm a_2275_11190# a_25054_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2773 a_23958_8154# row_n[6] a_24450_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2774 a_24962_15182# row_n[13] a_25454_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2775 a_8990_13174# a_2475_13198# a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2776 VDD rowon_n[7] a_6890_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2777 VDD rowon_n[15] a_7894_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2778 a_5374_14540# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2779 a_15414_14540# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2780 a_21950_3134# row_n[1] a_22442_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2781 a_9390_13536# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2782 a_2475_12194# a_1957_12194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X2783 a_5886_10162# row_n[8] a_6378_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2784 a_15926_10162# row_n[8] a_16418_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2785 a_26362_7190# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2786 a_27366_3174# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2787 a_33390_4178# rowon_n[2] a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2788 a_10998_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2789 a_17326_9198# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2790 a_27062_4138# a_2475_4162# a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2791 a_28978_6146# row_n[4] a_29470_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2792 a_24354_17230# rowon_n[15] a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2793 vcm a_2275_15206# a_13006_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2794 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2795 VSS row_n[1] a_12306_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2796 vcm a_2275_15206# a_2966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2797 a_32082_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2798 a_26970_1126# VDD a_27462_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2799 a_2161_18218# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2800 a_28370_16226# rowon_n[14] a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2801 VSS row_n[11] a_25358_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2802 a_22346_10202# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2803 a_2966_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2804 VDD rowon_n[2] a_32994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2805 a_14410_6508# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2806 a_20946_2130# a_2275_2154# a_21038_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2807 a_15318_12210# rowon_n[10] a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2808 a_16930_9158# row_n[7] a_17422_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2809 a_9294_8194# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2810 a_15014_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2811 a_31078_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2812 a_5278_12210# rowon_n[10] a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2813 VDD rowon_n[13] a_23958_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2814 a_12002_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2815 a_34090_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2816 a_21438_12532# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2817 a_10906_8154# a_2275_8178# a_10998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2818 a_18330_5182# rowon_n[3] a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2819 a_12402_1488# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2820 a_19334_1166# en_bit_n[2] a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2821 a_31382_1166# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2822 a_11910_4138# a_2275_4162# a_12002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2823 a_9294_11206# rowon_n[9] a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2824 VSS row_n[0] a_4274_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2825 a_30378_5182# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2826 a_25454_11528# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2827 VSS VDD a_17326_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2828 a_23350_18234# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2829 vcm a_2275_5166# a_34090_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2830 VDD rowon_n[8] a_14922_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2831 a_7986_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2832 VDD rowon_n[8] a_4882_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2833 a_6982_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2834 VSS row_n[15] a_3270_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2835 VSS row_n[15] a_13310_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2836 a_29982_3134# row_n[1] a_30474_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2837 VDD rowon_n[1] a_17934_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2838 VSS row_n[14] a_17326_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2839 a_22042_16186# a_2475_16210# a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2840 a_14314_13214# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2841 a_2874_7150# a_2275_7174# a_2966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2842 vcm a_2275_1150# a_9994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2843 a_3878_3134# a_2275_3158# a_3970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2844 VSS row_n[14] a_7286_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2845 a_13006_15182# a_2475_15206# a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2846 a_35094_15182# a_2475_15206# a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2847 a_4274_13214# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2848 vcm a_2275_12194# a_32082_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2849 a_23446_7512# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2850 a_15926_6146# a_2275_6170# a_16018_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2851 a_22954_16186# row_n[14] a_23446_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2852 a_2966_15182# a_2475_15206# a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2853 VSS row_n[7] a_27366_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2854 a_35398_3174# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2855 a_9902_14178# a_2275_14202# a_9994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2856 a_17022_14178# a_2475_14202# a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2857 a_21438_2492# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2858 VDD VDD a_15926_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2859 a_13406_15544# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2860 a_6982_14178# a_2475_14202# a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2861 VDD VDD a_5886_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2862 a_3366_15544# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2863 VSS row_n[0] a_26362_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2864 a_2161_3158# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2865 a_13918_11166# row_n[9] a_14410_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2866 a_3878_11166# row_n[9] a_4370_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2867 vcm a_2275_9182# a_20034_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2868 a_35002_1126# VDD a_35494_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2869 a_26058_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2870 a_30074_9158# a_2475_9182# a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2871 VSS row_n[6] a_16322_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2872 a_7894_5142# a_2275_5166# a_7986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2873 a_8898_1126# a_2275_1150# a_8990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2874 a_27462_9520# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2875 a_28466_5504# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2876 a_23350_12210# rowon_n[10] a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2877 a_20946_10162# a_2275_10186# a_21038_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2878 a_6378_8516# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2879 a_13006_6146# a_2475_6170# a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2880 a_11302_2170# rowon_n[0] a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2881 a_22042_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2882 a_22346_18234# VDD a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2883 vcm a_2275_16210# a_10998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2884 a_35398_17230# rowon_n[15] a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2885 VDD rowon_n[3] a_12914_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2886 VSS row_n[12] a_23350_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2887 a_8990_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2888 a_23958_17190# a_2275_17214# a_24050_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2889 a_19430_12532# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2890 VDD rowon_n[8] a_22954_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2891 VSS row_n[5] a_8290_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2892 a_27974_16186# a_2275_16210# a_28066_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2893 a_32082_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2894 a_22346_6186# rowon_n[4] a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2895 a_4974_5142# a_2475_5166# a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2896 a_5978_1126# a_2475_1150# a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2897 VDD rowon_n[14] a_21950_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2898 VDD rowon_n[13] a_35002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2899 a_10298_6186# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2900 a_18026_4138# a_2475_4162# a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2901 a_35398_12210# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2902 a_17022_8154# a_2475_8178# a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2903 VSS row_n[10] a_12306_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2904 vcm a_2275_6170# a_14010_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2905 a_34394_18234# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2906 VSS VDD a_11302_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2907 a_34490_14540# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2908 a_34090_10162# a_2475_10186# a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2909 a_12002_10162# a_2475_10186# a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2910 vcm a_2275_18218# a_29070_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2911 VDD rowon_n[12] a_10906_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2912 a_12306_14218# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2913 a_35002_10162# row_n[8] a_35494_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2914 VSS row_n[0] a_34394_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2915 a_3270_1166# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2916 a_9994_3134# a_2475_3158# a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2917 a_27366_4178# rowon_n[2] a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2918 a_10998_16186# a_2475_16210# a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2919 a_33086_16186# a_2475_16210# a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2920 a_19334_10202# rowon_n[8] a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2921 a_26362_8194# rowon_n[6] a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2922 a_8990_7150# a_2475_7174# a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2923 vcm a_2275_2154# a_28066_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2924 a_15318_4178# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2925 a_33998_16186# row_n[14] a_34490_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2926 a_12402_10524# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2927 vcm a_2275_1150# a_6982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2928 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2929 a_10298_17230# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2930 vcm a_2275_5166# a_5978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2931 a_11398_16548# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2932 vcm a_2275_8178# a_18026_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2933 vcm a_2275_4162# a_19030_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2934 a_20034_4138# a_2475_4162# a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2935 a_26058_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2936 a_15318_7190# rowon_n[5] a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2937 a_32994_7150# a_2275_7174# a_33086_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2938 a_33998_3134# a_2275_3158# a_34090_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2939 a_21950_6146# row_n[4] a_22442_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2940 VDD rowon_n[2] a_26970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2941 a_2475_15206# a_1957_15206# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X2942 VDD rowon_n[5] a_4882_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2943 a_14922_4138# row_n[2] a_15414_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2944 a_9902_15182# row_n[13] a_10394_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2945 a_21342_13214# rowon_n[11] a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2946 vcm a_2275_11190# a_9994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2947 a_34394_12210# rowon_n[10] a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2948 a_31990_10162# a_2275_10186# a_32082_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2949 a_9294_9198# rowon_n[7] a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2950 a_22954_12170# a_2275_12194# a_23046_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2951 a_24354_5182# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2952 a_24050_6146# a_2475_6170# a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2953 a_21950_18194# a_2275_18218# a_22042_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2954 VDD rowon_n[9] a_20946_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2955 VDD rowon_n[8] a_33998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2956 a_25966_8154# row_n[6] a_26458_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2957 VDD rowon_n[7] a_8898_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2958 VSS VDD a_10298_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2959 VSS row_n[15] a_32386_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2960 a_23958_3134# row_n[1] a_24450_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2961 a_20338_14218# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2962 a_2475_16210# a_1957_16210# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X2963 a_33390_13214# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2964 a_12002_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2965 a_28370_7190# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2966 a_29374_3174# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2967 a_13006_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2968 a_27062_17190# a_2475_17214# a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2969 a_3270_16226# rowon_n[14] a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2970 a_13310_16226# rowon_n[14] a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2971 VSS row_n[11] a_10298_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2972 a_7286_6186# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2973 a_29070_4138# a_2475_4162# a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2974 a_19334_9198# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2975 a_27974_17190# row_n[15] a_28466_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2976 a_32482_15544# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2977 vcm a_2275_13198# a_28066_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2978 a_32082_11166# a_2475_11190# a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2979 a_4882_15182# a_2275_15206# a_4974_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2980 a_14922_15182# a_2275_15206# a_15014_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2981 VSS row_n[7] a_20338_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2982 a_30378_9198# rowon_n[7] a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2983 VSS row_n[1] a_14314_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2984 a_32994_11166# row_n[9] a_33486_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2985 a_28978_1126# VDD a_29470_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2986 vcm a_2275_3158# a_32082_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2987 a_10394_11528# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2988 a_34090_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2989 vcm a_2275_7174# a_31078_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2990 VDD rowon_n[4] a_17934_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2991 a_29982_6146# row_n[4] a_30474_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2992 a_8898_12170# row_n[10] a_9390_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2993 a_18938_12170# row_n[10] a_19430_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2994 a_3970_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2995 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2996 a_4974_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2997 a_17022_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2998 a_22954_2130# a_2275_2154# a_23046_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2999 VDD a_2161_4162# a_2275_4162# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X3000 a_2161_13198# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3001 a_18938_9158# row_n[7] a_19430_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3002 a_33086_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3003 vcm a_2275_16210# a_30074_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3004 a_20434_9520# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3005 a_12914_8154# a_2275_8178# a_13006_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3006 a_14410_1488# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3007 a_13918_4138# a_2275_4162# a_14010_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3008 a_21438_5504# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3009 VDD rowon_n[7] a_29982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3010 a_33390_1166# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3011 vcm a_2275_17214# a_16018_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3012 vcm a_2275_17214# a_5978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3013 VSS row_n[13] a_28370_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3014 a_32386_13214# rowon_n[11] a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3015 a_20034_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3016 a_8990_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3017 a_9994_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3018 a_29374_11206# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3019 a_24050_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3020 a_20946_13174# a_2275_13198# a_21038_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3021 a_4882_7150# a_2275_7174# a_4974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3022 a_5886_3134# a_2275_3158# a_5978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3023 VDD rowon_n[15] a_26970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3024 a_15014_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3025 a_33998_12170# a_2275_12194# a_34090_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3026 a_25454_7512# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3027 a_17934_6146# a_2275_6170# a_18026_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3028 a_4974_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3029 VDD rowon_n[5] a_35002_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3030 a_8990_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3031 a_28466_13536# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3032 VDD rowon_n[9] a_31990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3033 VSS row_n[7] a_29374_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3034 a_10998_4138# a_2475_4162# a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3035 a_23446_2492# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3036 VSS VDD a_30378_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3037 VSS row_n[0] a_28370_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3038 a_31382_14218# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3039 a_32386_8194# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3040 VSS row_n[3] a_6282_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3041 a_1957_2154# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3042 a_25054_18194# a_2475_18218# a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3043 vcm a_2275_15206# a_22042_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3044 a_32082_9158# a_2475_9182# a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3045 VSS row_n[6] a_18330_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3046 a_16018_17190# a_2475_17214# a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3047 a_7286_15222# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3048 a_17326_15222# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3049 a_29470_9520# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3050 a_25966_18194# VDD a_26458_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3051 a_5978_17190# a_2475_17214# a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3052 vcm a_2275_14202# a_26058_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3053 a_8386_8516# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3054 a_2966_3134# a_2475_3158# a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3055 a_20338_4178# rowon_n[2] a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3056 a_12914_16186# a_2275_16210# a_13006_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3057 a_30474_16548# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3058 a_15014_6146# a_2475_6170# a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3059 vcm a_2275_2154# a_21038_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3060 a_13310_2170# rowon_n[0] a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3061 a_24050_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3062 a_2874_16186# a_2275_16210# a_2966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3063 a_9994_16186# a_2475_16210# a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3064 a_26970_7150# a_2275_7174# a_27062_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3065 a_31078_2130# a_2475_2154# a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3066 a_6378_17552# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3067 a_16418_17552# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3068 vcm a_2275_8178# a_10998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3069 a_6378_3496# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3070 vcm a_2275_4162# a_12002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3071 a_16930_13174# row_n[11] a_17422_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3072 a_6890_13174# row_n[11] a_7382_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3073 VDD rowon_n[2] a_19942_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3074 vcm a_2275_12194# a_15014_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3075 vcm a_2275_12194# a_4974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3076 a_24354_6186# rowon_n[4] a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3077 a_6982_5142# a_2475_5166# a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3078 a_7986_1126# a_2475_1150# a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3079 VSS row_n[8] a_27366_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3080 vcm a_2275_18218# a_3970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3081 vcm a_2275_18218# a_14010_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3082 a_27974_11166# a_2275_11190# a_28066_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3083 vcm a_2275_7174# a_2966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3084 vcm a_2275_3158# a_3970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3085 vcm a_2275_6170# a_16018_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3086 VSS row_n[14] a_26362_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3087 a_30378_14218# rowon_n[12] a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3088 VDD rowon_n[10] a_25966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3089 a_31990_1126# a_2275_1150# a_32082_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3090 a_30986_5142# a_2275_5166# a_31078_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3091 a_31078_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3092 a_35094_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3093 a_31990_13174# a_2275_13198# a_32082_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3094 a_5278_1166# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3095 VSS row_n[2] a_19334_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3096 VDD VDD a_24962_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3097 a_2966_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3098 a_13006_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3099 a_28370_8194# rowon_n[6] a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3100 a_29374_4178# rowon_n[2] a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3101 a_25358_15222# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3102 VDD rowon_n[6] a_14922_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3103 vcm a_2275_5166# a_7986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3104 vcm a_2275_1150# a_8990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3105 a_21342_7190# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3106 a_22346_3174# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3107 a_8290_17230# rowon_n[15] a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3108 VDD a_2161_11190# a_2275_11190# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X3109 VSS row_n[5] a_31382_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3110 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=2.7645 pd=21.91 as=0.2755 ps=2.19 w=1.9 l=0.22 M=2
X3111 a_24450_17552# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3112 a_20946_14178# row_n[12] a_21438_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3113 VSS row_n[11] a_9294_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3114 a_24050_13174# a_2475_13198# a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3115 a_6282_10202# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3116 a_16322_10202# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3117 vcm a_2275_10186# a_21038_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3118 a_12306_9198# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3119 a_35002_7150# a_2275_7174# a_35094_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3120 a_22042_4138# a_2475_4162# a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3121 a_4974_12170# a_2475_12194# a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3122 a_15014_12170# a_2475_12194# a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3123 a_28066_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3124 a_17326_7190# rowon_n[5] a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3125 a_23958_6146# row_n[4] a_24450_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3126 VDD rowon_n[2] a_28978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3127 a_19430_4500# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3128 a_24962_13174# row_n[11] a_25454_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3129 a_8990_11166# a_2475_11190# a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3130 VDD rowon_n[5] a_6890_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3131 VDD rowon_n[13] a_7894_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3132 a_5374_12532# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3133 a_15414_12532# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3134 a_21950_1126# VDD a_22442_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3135 VDD rowon_n[0] a_4882_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3136 a_9390_11528# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3137 a_2475_10186# a_1957_10186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X3138 a_27366_1166# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3139 a_26362_5182# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3140 a_11910_9158# row_n[7] a_12402_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3141 a_4274_8194# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3142 vcm a_2275_17214# a_35094_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3143 a_27974_8154# row_n[6] a_28466_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3144 a_12914_17190# row_n[15] a_13406_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3145 a_24354_15222# rowon_n[13] a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3146 vcm a_2275_13198# a_13006_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3147 VSS row_n[10] a_21342_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3148 VSS VDD a_12306_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3149 a_2874_17190# row_n[15] a_3366_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3150 vcm a_2275_13198# a_2966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3151 a_25966_3134# row_n[1] a_26458_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3152 a_28370_14218# rowon_n[12] a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3153 VSS row_n[9] a_25358_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3154 a_2966_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3155 a_15014_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3156 a_29070_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3157 VDD rowon_n[12] a_19942_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3158 a_30074_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3159 a_15318_10202# rowon_n[8] a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3160 a_14010_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3161 a_16930_7150# row_n[5] a_17422_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3162 a_9294_6186# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3163 a_5278_10202# rowon_n[8] a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3164 VDD rowon_n[11] a_23958_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3165 a_21438_10524# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3166 a_10906_6146# a_2275_6170# a_10998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3167 a_18330_3174# rowon_n[1] a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3168 VSS row_n[7] a_22346_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3169 a_30378_3174# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3170 a_32386_9198# rowon_n[7] a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3171 a_23350_16226# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3172 vcm a_2275_7174# a_33086_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3173 vcm a_2275_3158# a_34090_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3174 a_14922_10162# a_2275_10186# a_15014_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3175 a_26058_9158# a_2475_9182# a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3176 VSS row_n[0] a_21342_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3177 a_6982_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3178 a_4882_10162# a_2275_10186# a_4974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3179 a_6282_18234# VDD a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3180 a_16322_18234# VDD a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3181 VSS row_n[13] a_3270_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3182 VSS row_n[13] a_13310_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3183 a_35094_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3184 a_3878_1126# a_2275_1150# a_3970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3185 VDD en_bit_n[1] a_17934_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3186 a_29982_1126# VDD a_30474_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3187 a_24962_2130# a_2275_2154# a_25054_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3188 a_22442_18556# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3189 VSS row_n[12] a_17326_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3190 a_22042_14178# a_2475_14202# a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3191 a_14314_11206# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3192 VSS row_n[6] a_11302_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3193 a_2874_5142# a_2275_5166# a_2966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3194 a_35494_17552# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3195 VSS row_n[12] a_7286_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3196 a_31990_14178# row_n[12] a_32482_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3197 a_13006_13174# a_2475_13198# a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3198 a_35094_13174# a_2475_13198# a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3199 a_4274_11206# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3200 vcm a_2275_10186# a_32082_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3201 a_22442_9520# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3202 a_14922_8154# a_2275_8178# a_15014_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3203 a_35398_1166# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15 M=2
X3204 a_15926_4138# a_2275_4162# a_16018_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3205 a_23446_5504# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3206 a_17934_17190# a_2275_17214# a_18026_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3207 a_2966_13174# a_2475_13198# a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3208 VDD rowon_n[7] a_31990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3209 a_7894_17190# a_2275_17214# a_7986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3210 VDD rowon_n[15] a_11910_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3211 VDD rowon_n[14] a_15926_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3212 a_13406_13536# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3213 VDD rowon_n[14] a_5886_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3214 a_3366_13536# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3215 VSS row_n[5] a_3270_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3216 vcm a_2275_18218# a_33086_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3217 VSS row_n[4] a_16322_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3218 a_7894_3134# a_2275_3158# a_7986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3219 VSS row_n[10] a_19334_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3220 a_27462_7512# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3221 a_24050_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3222 a_23350_10202# rowon_n[8] a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3223 a_6378_6508# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3224 a_13006_4138# a_2475_4162# a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3225 a_15014_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3226 a_12002_8154# a_2475_8178# a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3227 a_25454_2492# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3228 a_10906_18194# VDD a_11398_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3229 a_22346_16226# rowon_n[14] a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3230 a_35398_15222# rowon_n[13] a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3231 vcm a_2275_14202# a_10998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3232 a_4974_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3233 VDD rowon_n[0] a_35002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3234 VDD rowon_n[12] a_17934_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3235 a_34394_8194# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3236 a_27062_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3237 a_23958_15182# a_2275_15206# a_24050_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3238 a_19430_10524# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3239 VSS row_n[3] a_8290_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3240 a_18026_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3241 a_34090_9158# a_2475_9182# a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3242 a_7986_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3243 a_27974_14178# a_2275_14202# a_28066_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3244 a_21342_8194# rowon_n[6] a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3245 a_4974_3134# a_2475_3158# a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3246 a_22346_4178# rowon_n[2] a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3247 VDD rowon_n[11] a_35002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3248 a_3970_7150# a_2475_7174# a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3249 vcm a_2275_2154# a_23046_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3250 a_10298_4178# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3251 a_35398_10202# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3252 a_17022_6146# a_2475_6170# a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3253 a_33086_2130# a_2475_2154# a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3254 a_28978_7150# a_2275_7174# a_29070_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3255 a_8386_3496# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3256 VSS row_n[8] a_12306_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3257 vcm a_2275_8178# a_13006_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3258 vcm a_2275_4162# a_14010_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3259 a_34394_16226# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3260 a_2874_11166# a_2275_11190# a_2966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3261 a_12914_11166# a_2275_11190# a_13006_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3262 VSS row_n[14] a_11302_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3263 a_34490_12532# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3264 a_21038_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3265 a_10298_7190# rowon_n[5] a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3266 VDD rowon_n[2] a_21950_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3267 vcm a_2275_16210# a_29070_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3268 a_33086_14178# a_2475_14202# a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3269 VDD rowon_n[10] a_10906_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3270 a_26362_6186# rowon_n[4] a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3271 a_9994_1126# a_2475_1150# a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3272 a_9902_4138# row_n[2] a_10394_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3273 a_33486_18556# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3274 a_10998_14178# a_2475_14202# a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3275 a_8990_5142# a_2475_5166# a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3276 a_5886_18194# a_2275_18218# a_5978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3277 VDD VDD a_9902_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3278 a_15926_18194# a_2275_18218# a_16018_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3279 a_4274_9198# rowon_n[7] a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3280 a_10298_15222# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3281 vcm a_2275_7174# a_4974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3282 vcm a_2275_3158# a_5978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3283 vcm a_2275_6170# a_18026_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3284 a_2475_2154# a_1957_2154# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X3285 a_15318_5182# rowon_n[3] a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3286 a_32994_5142# a_2275_5166# a_33086_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3287 a_20946_8154# row_n[6] a_21438_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3288 VDD rowon_n[7] a_3878_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3289 a_31478_8516# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3290 VDD rowon_n[3] a_4882_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3291 a_9902_13174# row_n[11] a_10394_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3292 a_21342_11206# rowon_n[9] a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3293 VDD rowon_n[6] a_16930_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3294 a_35094_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3295 a_34394_10202# rowon_n[8] a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3296 a_2966_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3297 a_13006_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3298 a_23350_7190# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3299 a_24354_3174# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3300 VDD rowon_n[1] a_14922_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3301 VDD rowon_n[12] a_28978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3302 a_17022_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3303 VSS row_n[5] a_33390_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3304 a_24050_4138# a_2475_4162# a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3305 a_6982_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3306 a_14314_9198# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3307 vcm a_2275_7174# a_27062_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3308 a_21950_16186# a_2275_16210# a_22042_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3309 a_25966_6146# row_n[4] a_26458_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3310 a_5978_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3311 a_16018_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3312 VDD rowon_n[5] a_8898_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3313 a_28370_17230# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3314 VSS row_n[13] a_32386_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3315 a_23958_1126# VDD a_24450_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3316 a_2475_14202# a_1957_14202# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X3317 a_33390_11206# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3318 VDD rowon_n[0] a_6890_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3319 a_13310_14218# rowon_n[12] a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3320 a_12002_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3321 a_29374_1166# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3322 a_28370_5182# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3323 VDD rowon_n[15] a_30986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3324 a_27062_15182# a_2475_15206# a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3325 a_3270_14218# rowon_n[12] a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3326 a_9294_12210# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3327 a_19334_12210# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3328 vcm a_2275_12194# a_24050_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3329 VSS row_n[9] a_10298_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3330 a_13918_9158# row_n[7] a_14410_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3331 a_6282_8194# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3332 a_7286_4178# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3333 vcm a_2275_11190# a_28066_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3334 a_27974_15182# row_n[13] a_28466_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3335 a_32482_13536# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3336 a_4882_13174# a_2275_13198# a_4974_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3337 a_14922_13174# a_2275_13198# a_15014_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3338 VSS VDD a_14314_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3339 a_8386_14540# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3340 a_18426_14540# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3341 vcm a_2275_1150# a_32082_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3342 a_27974_3134# row_n[1] a_28466_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3343 vcm a_2275_5166# a_31078_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3344 a_8898_10162# row_n[8] a_9390_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3345 a_18938_10162# row_n[8] a_19430_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3346 a_3970_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3347 a_4974_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3348 a_6890_4138# row_n[2] a_7382_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3349 a_17022_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3350 a_18938_7150# row_n[5] a_19430_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3351 a_29982_18194# VDD a_30474_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3352 vcm a_2275_14202# a_30074_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3353 a_20434_7512# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3354 a_12914_6146# a_2275_6170# a_13006_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3355 VDD rowon_n[5] a_29982_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3356 a_16930_2130# row_n[0] a_17422_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3357 a_27366_17230# rowon_n[15] a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3358 vcm a_2275_15206# a_16018_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3359 VSS row_n[7] a_24354_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3360 vcm a_2275_15206# a_5978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3361 a_34394_9198# rowon_n[7] a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3362 VSS row_n[11] a_28370_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3363 a_32386_11206# rowon_n[9] a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3364 a_28066_9158# a_2475_9182# a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3365 vcm a_2275_7174# a_35094_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3366 a_20034_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3367 VSS row_n[0] a_23350_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3368 a_8990_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3369 a_24050_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3370 VSS row_n[6] a_13310_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3371 a_19030_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3372 a_4882_5142# a_2275_5166# a_4974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3373 a_5886_1126# a_2275_1150# a_5978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3374 VDD rowon_n[13] a_26970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3375 a_15014_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3376 a_24450_9520# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3377 a_17934_4138# a_2275_4162# a_18026_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3378 a_25454_5504# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3379 a_4974_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3380 VDD rowon_n[7] a_33998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3381 a_3366_8516# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3382 VDD rowon_n[3] a_35002_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3383 a_28466_11528# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3384 VSS a_2161_9182# a_2275_9182# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X3385 a_21950_7150# a_2275_7174# a_22042_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3386 a_26362_18234# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3387 VSS row_n[14] a_30378_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3388 VSS row_n[15] a_6282_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3389 VSS row_n[15] a_16322_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3390 a_21038_17190# a_2475_17214# a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3391 VSS row_n[5] a_5278_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3392 a_32386_6186# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3393 VSS row_n[1] a_6282_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3394 a_35002_18194# a_2275_18218# a_35094_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3395 a_25054_16186# a_2475_16210# a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3396 a_17326_13214# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3397 vcm a_2275_13198# a_22042_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3398 VSS row_n[4] a_18330_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3399 a_21950_17190# row_n[15] a_22442_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3400 a_1957_16210# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3401 a_16018_15182# a_2475_15206# a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3402 a_7286_13214# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3403 a_29470_7512# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3404 a_25966_16186# row_n[14] a_26458_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3405 a_5978_15182# a_2475_15206# a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3406 a_8386_6508# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3407 a_2966_1126# a_2475_1150# a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3408 a_12914_14178# a_2275_14202# a_13006_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3409 a_14010_8154# a_2475_8178# a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3410 a_15014_4138# a_2475_4162# a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3411 a_16418_15544# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3412 a_2874_14178# a_2275_14202# a_2966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3413 a_9994_14178# a_2475_14202# a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3414 a_27462_2492# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3415 a_26970_5142# a_2275_5166# a_27062_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3416 VDD VDD a_8898_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3417 a_6378_15544# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3418 vcm a_2275_6170# a_10998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3419 a_6378_1488# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3420 a_16930_11166# row_n[9] a_17422_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3421 a_6890_11166# row_n[9] a_7382_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3422 vcm a_2275_10186# a_15014_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3423 a_4882_14178# row_n[12] a_5374_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3424 a_14922_14178# row_n[12] a_15414_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3425 a_26362_12210# rowon_n[10] a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3426 vcm a_2275_10186# a_4974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3427 a_23958_10162# a_2275_10186# a_24050_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3428 a_23350_8194# rowon_n[6] a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3429 a_6982_3134# a_2475_3158# a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3430 a_24354_4178# rowon_n[2] a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3431 VDD rowon_n[6] a_9902_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3432 vcm a_2275_2154# a_25054_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3433 a_25358_18234# VDD a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3434 a_1957_17214# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3435 vcm a_2275_16210# a_3970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3436 vcm a_2275_16210# a_14010_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3437 vcm a_2275_5166# a_2966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3438 a_35094_2130# a_2475_2154# a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3439 vcm a_2275_1150# a_3970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3440 vcm a_2275_8178# a_15014_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3441 vcm a_2275_4162# a_16018_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3442 VSS row_n[12] a_26362_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3443 a_26970_17190# a_2275_17214# a_27062_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3444 VDD rowon_n[8] a_25966_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3445 a_29982_7150# a_2275_7174# a_30074_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3446 a_30986_3134# a_2275_3158# a_31078_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3447 a_31078_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3448 a_23046_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3449 a_12306_7190# rowon_n[5] a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3450 VDD rowon_n[2] a_23958_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3451 VSS row_n[15] a_24354_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3452 a_35094_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3453 VDD rowon_n[14] a_24962_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3454 a_2966_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3455 a_13006_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3456 a_28370_6186# rowon_n[4] a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3457 a_25358_13214# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3458 a_6282_9198# rowon_n[7] a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3459 VDD rowon_n[4] a_14922_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3460 vcm a_2275_3158# a_7986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3461 a_19030_17190# a_2475_17214# a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3462 VSS row_n[10] a_15318_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3463 a_20034_12170# a_2475_12194# a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3464 a_22346_1166# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3465 a_21342_5182# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3466 a_8290_15222# rowon_n[13] a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3467 VSS row_n[10] a_5278_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3468 a_5278_2170# rowon_n[0] a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3469 VSS row_n[3] a_31382_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3470 a_24450_15544# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3471 a_20946_12170# row_n[10] a_21438_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3472 VSS row_n[9] a_9294_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3473 a_24050_11166# a_2475_11190# a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3474 a_35002_5142# a_2275_5166# a_35094_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3475 a_4974_10162# a_2475_10186# a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3476 a_15014_10162# a_2475_10186# a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3477 a_22954_8154# row_n[6] a_23446_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3478 a_17326_5182# rowon_n[3] a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3479 VDD rowon_n[12] a_13918_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3480 a_24962_11166# row_n[9] a_25454_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3481 a_33486_8516# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3482 VDD rowon_n[12] a_3878_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3483 VDD rowon_n[7] a_5886_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3484 VDD rowon_n[3] a_6890_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3485 VDD rowon_n[11] a_7894_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3486 a_5374_10524# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3487 a_15414_10524# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3488 a_20946_3134# row_n[1] a_21438_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3489 a_13310_17230# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3490 a_31478_3496# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3491 a_3270_17230# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3492 a_26362_3174# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3493 VDD rowon_n[1] a_16930_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3494 a_11910_7150# row_n[5] a_12402_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3495 a_25358_7190# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3496 VSS row_n[5] a_35398_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3497 a_4274_6186# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3498 vcm a_2275_15206# a_35094_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3499 a_16322_9198# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3500 vcm a_2275_7174# a_29070_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3501 a_27974_6146# row_n[4] a_28466_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3502 a_12914_15182# row_n[13] a_13406_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3503 a_24354_13214# rowon_n[11] a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3504 vcm a_2275_11190# a_13006_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3505 VSS row_n[8] a_21342_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3506 a_2874_15182# row_n[13] a_3366_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3507 vcm a_2275_11190# a_2966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3508 a_21950_11166# a_2275_11190# a_22042_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3509 a_25966_1126# VDD a_26458_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3510 a_21038_9158# a_2475_9182# a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3511 VDD rowon_n[0] a_8898_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3512 VDD rowon_n[15] a_18938_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3513 a_29070_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3514 VDD rowon_n[10] a_19942_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3515 a_25966_12170# a_2275_12194# a_26058_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3516 a_15926_9158# row_n[7] a_16418_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3517 a_14010_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3518 a_16930_5142# row_n[3] a_17422_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3519 a_30074_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3520 a_19942_2130# a_2275_2154# a_20034_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3521 a_9294_4178# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3522 a_8290_8194# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3523 VDD rowon_n[9] a_23958_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3524 a_9902_8154# a_2275_8178# a_9994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3525 a_18330_1166# en_bit_n[1] a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3526 a_30378_1166# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3527 a_10906_4138# a_2275_4162# a_10998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3528 VSS VDD a_22346_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3529 VSS row_n[15] a_35398_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3530 a_23350_14218# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3531 vcm a_2275_5166# a_33086_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3532 a_12306_17230# rowon_n[15] a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3533 a_6982_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3534 a_8898_4138# row_n[2] a_9390_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3535 a_6282_16226# rowon_n[14] a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3536 a_16322_16226# rowon_n[14] a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3537 VSS row_n[11] a_3270_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3538 VSS row_n[11] a_13310_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3539 a_31078_12170# a_2475_12194# a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3540 a_22442_16548# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3541 VSS row_n[4] a_11302_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3542 a_2874_3134# a_2275_3158# a_2966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3543 a_35494_15544# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3544 a_31990_12170# row_n[10] a_32482_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3545 a_13006_11166# a_2475_11190# a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3546 a_35094_11166# a_2475_11190# a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3547 a_22442_7512# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3548 a_14922_6146# a_2275_6170# a_15014_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3549 a_7894_15182# a_2275_15206# a_7986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3550 a_17934_15182# a_2275_15206# a_18026_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3551 a_2966_11166# a_2475_11190# a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3552 VDD rowon_n[5] a_31990_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3553 a_18938_2130# row_n[0] a_19430_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3554 VDD rowon_n[13] a_11910_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3555 a_20434_2492# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3556 a_13406_11528# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3557 VDD rowon_n[0] a_29982_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3558 a_3366_11528# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3559 a_11302_18234# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3560 a_35398_2170# rowon_n[0] a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3561 VSS row_n[0] a_25358_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3562 VSS row_n[3] a_3270_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3563 vcm a_2275_16210# a_33086_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3564 a_20034_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3565 VSS row_n[6] a_15318_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3566 a_7894_1126# a_2275_1150# a_7986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3567 VSS row_n[2] a_16322_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3568 VSS row_n[8] a_19334_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3569 a_27462_5504# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3570 vcm a_2275_17214# a_19030_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3571 a_5374_8516# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3572 a_5978_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3573 vcm a_2275_17214# a_8990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3574 a_12002_6146# a_2475_6170# a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3575 a_10906_16186# row_n[14] a_11398_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3576 a_22346_14218# rowon_n[12] a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3577 a_35398_13214# rowon_n[11] a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3578 a_23958_7150# a_2275_7174# a_24050_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3579 a_3366_3496# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3580 a_23046_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3581 VDD rowon_n[10] a_17934_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3582 a_34394_6186# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3583 a_16418_4500# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3584 a_27062_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3585 a_23958_13174# a_2275_13198# a_24050_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3586 VSS row_n[5] a_7286_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3587 VSS row_n[1] a_8290_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3588 a_18026_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3589 a_1957_8178# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3590 a_7986_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3591 a_21342_6186# rowon_n[4] a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3592 a_4974_1126# a_2475_1150# a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3593 a_2161_2154# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3594 VSS row_n[10] a_34394_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3595 VDD rowon_n[9] a_35002_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3596 a_3970_5142# a_2475_5166# a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3597 a_11302_12210# rowon_n[10] a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3598 a_1957_11190# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3599 a_17022_4138# a_2475_4162# a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3600 VSS VDD a_33390_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3601 a_8386_1488# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3602 a_29470_2492# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3603 a_28978_5142# a_2275_5166# a_29070_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3604 a_29070_12170# a_2475_12194# a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3605 a_6890_8154# a_2275_8178# a_6982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3606 vcm a_2275_6170# a_13006_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3607 a_10298_18234# VDD a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3608 VDD rowon_n[12] a_32994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3609 a_34394_14218# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3610 a_28066_18194# a_2475_18218# a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3611 VSS row_n[12] a_11302_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3612 a_34490_10524# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3613 a_10298_5182# rowon_n[3] a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3614 a_28978_18194# VDD a_29470_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3615 a_11910_17190# a_2275_17214# a_12002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3616 vcm a_2275_14202# a_29070_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3617 VDD rowon_n[8] a_10906_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3618 a_26362_4178# rowon_n[2] a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3619 a_15926_16186# a_2275_16210# a_16018_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3620 a_33486_16548# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3621 VDD rowon_n[6] a_11910_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3622 a_8990_3134# a_2475_3158# a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3623 a_5886_16186# a_2275_16210# a_5978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3624 VDD rowon_n[14] a_9902_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3625 a_19030_8154# a_2475_8178# a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3626 a_10298_13214# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3627 vcm a_2275_5166# a_4974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3628 vcm a_2275_1150# a_5978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3629 VDD rowon_n[1] a_9902_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3630 vcm a_2275_4162# a_18026_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3631 a_25054_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3632 a_14314_7190# rowon_n[5] a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3633 vcm a_2275_7174# a_22042_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3634 a_32994_3134# a_2275_3158# a_33086_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3635 a_15318_3174# rowon_n[1] a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3636 vcm a_2275_12194# a_18026_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3637 a_20946_6146# row_n[4] a_21438_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3638 VDD rowon_n[2] a_25966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3639 vcm a_2275_12194# a_7986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3640 VDD rowon_n[5] a_3878_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3641 a_31478_6508# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3642 a_9902_11166# row_n[9] a_10394_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3643 a_31078_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3644 VDD rowon_n[4] a_16930_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3645 vcm a_2275_18218# a_6982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3646 vcm a_2275_18218# a_17022_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3647 a_8290_9198# rowon_n[7] a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3648 a_22042_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3649 VDD VSS a_14922_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3650 a_24354_1166# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3651 a_23350_5182# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3652 a_21038_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3653 VDD rowon_n[10] a_28978_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3654 a_7286_2170# rowon_n[0] a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3655 VSS row_n[3] a_33390_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3656 vcm a_2275_5166# a_27062_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3657 a_31382_17230# rowon_n[15] a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3658 a_21950_14178# a_2275_14202# a_22042_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3659 a_24962_8154# row_n[6] a_25454_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3660 a_5978_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3661 a_16018_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3662 VDD rowon_n[7] a_7894_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3663 a_35494_8516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3664 VDD rowon_n[3] a_8898_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3665 a_28370_15222# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3666 VSS row_n[11] a_32386_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3667 a_19942_17190# a_2275_17214# a_20034_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3668 a_33486_3496# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3669 a_22954_3134# row_n[1] a_23446_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3670 a_28370_3174# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3671 a_12002_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3672 a_27462_17552# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3673 VDD rowon_n[13] a_30986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3674 a_23958_14178# row_n[12] a_24450_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3675 a_27062_13174# a_2475_13198# a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3676 a_9294_10202# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3677 a_19334_10202# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3678 vcm a_2275_10186# a_24050_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3679 a_13918_7150# row_n[5] a_14410_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3680 a_6282_6186# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3681 a_7986_12170# a_2475_12194# a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3682 a_10906_12170# a_2275_12194# a_10998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3683 a_18026_12170# a_2475_12194# a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3684 a_18330_9198# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3685 a_27974_13174# row_n[11] a_28466_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3686 a_32482_11528# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3687 a_11910_2130# row_n[0] a_12402_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3688 a_30378_18234# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3689 a_8386_12532# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3690 a_18426_12532# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3691 a_17326_2170# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3692 a_23046_9158# a_2475_9182# a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3693 vcm a_2275_7174# a_30074_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3694 a_27974_1126# VDD a_28466_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3695 vcm a_2275_3158# a_31078_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3696 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3697 a_3970_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3698 vcm a_2275_18218# a_25054_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3699 a_17934_9158# row_n[7] a_18426_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3700 a_18938_5142# row_n[3] a_19430_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3701 a_32082_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3702 a_29982_16186# row_n[14] a_30474_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3703 a_12914_4138# a_2275_4162# a_13006_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3704 a_20434_5504# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3705 a_29070_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3706 VDD rowon_n[3] a_29982_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3707 a_15926_17190# row_n[15] a_16418_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3708 a_27366_15222# rowon_n[13] a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3709 vcm a_2275_13198# a_16018_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3710 a_5886_17190# row_n[15] a_6378_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3711 vcm a_2275_13198# a_5978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3712 VSS row_n[9] a_28370_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3713 vcm a_2275_5166# a_35094_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3714 a_19030_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3715 a_20034_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3716 a_8990_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3717 a_10998_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3718 a_33086_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3719 VSS row_n[4] a_13310_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3720 a_19030_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3721 a_4882_3134# a_2275_3158# a_4974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3722 VDD rowon_n[11] a_26970_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3723 a_24450_7512# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3724 VDD rowon_n[5] a_33998_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3725 a_3366_6508# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3726 a_22346_17230# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3727 a_2161_12194# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3728 a_16018_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3729 VSS a_2161_7174# a_2275_7174# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X3730 a_22442_2492# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3731 a_21950_5142# a_2275_5166# a_22042_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3732 a_26362_16226# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3733 VSS row_n[12] a_30378_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3734 a_17934_10162# a_2275_10186# a_18026_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3735 VDD rowon_n[0] a_31990_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3736 a_30986_17190# a_2275_17214# a_31078_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3737 a_7894_10162# a_2275_10186# a_7986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3738 VSS row_n[0] a_27366_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3739 a_9294_18234# VDD a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3740 VSS row_n[13] a_6282_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3741 VSS row_n[13] a_16322_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3742 a_21038_15182# a_2475_15206# a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3743 a_19334_8194# rowon_n[6] a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3744 a_31382_8194# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3745 VSS row_n[3] a_5278_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3746 VSS VDD a_6282_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3747 a_32386_4178# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3748 a_35002_16186# a_2275_16210# a_35094_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3749 a_25054_14178# a_2475_14202# a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3750 a_17326_11206# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3751 vcm a_2275_11190# a_22042_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3752 VSS row_n[2] a_18330_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3753 a_25454_18556# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3754 a_21950_15182# row_n[13] a_22442_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3755 a_1957_14202# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3756 a_16018_13174# a_2475_13198# a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3757 a_7286_11206# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3758 VSS row_n[6] a_17326_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3759 a_29470_5504# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3760 a_5978_13174# a_2475_13198# a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3761 a_7382_8516# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3762 VDD rowon_n[15] a_4882_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3763 VDD rowon_n[15] a_14922_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3764 a_7986_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3765 a_14010_6146# a_2475_6170# a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3766 vcm a_2275_2154# a_20034_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3767 a_16418_13536# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3768 a_25966_7150# a_2275_7174# a_26058_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3769 a_30074_2130# a_2475_2154# a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3770 a_26970_3134# a_2275_3158# a_27062_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3771 VDD rowon_n[14] a_8898_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3772 a_6378_13536# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3773 vcm a_2275_8178# a_9994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3774 a_5374_3496# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3775 a_31990_4138# row_n[2] a_32482_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3776 vcm a_2275_4162# a_10998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3777 a_16930_9158# a_2275_9182# a_17022_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3778 a_18426_4500# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3779 VSS row_n[5] a_9294_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3780 a_4882_12170# row_n[10] a_5374_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3781 a_14922_12170# row_n[10] a_15414_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3782 a_27062_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3783 a_26362_10202# rowon_n[8] a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3784 a_23350_6186# rowon_n[4] a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3785 a_6982_1126# a_2475_1150# a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3786 a_18026_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3787 VDD rowon_n[4] a_9902_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3788 a_3878_18194# VDD a_4370_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3789 a_13918_18194# VDD a_14410_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3790 a_25358_16226# rowon_n[14] a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3791 a_1957_15206# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3792 vcm a_2275_14202# a_3970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3793 vcm a_2275_14202# a_14010_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3794 a_7986_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3795 vcm a_2275_3158# a_2966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3796 a_8898_8154# a_2275_8178# a_8990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3797 vcm a_2275_6170# a_15014_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3798 a_26970_15182# a_2275_15206# a_27062_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3799 a_31078_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3800 a_30986_1126# a_2275_1150# a_31078_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3801 a_29982_5142# a_2275_5166# a_30074_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3802 a_12306_5182# rowon_n[3] a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3803 VSS row_n[13] a_24354_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3804 a_21342_12210# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3805 a_28370_4178# rowon_n[2] a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3806 a_25358_11206# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3807 VDD rowon_n[6] a_13918_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3808 vcm a_2275_1150# a_7986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3809 VDD rowon_n[15] a_22954_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3810 a_19030_15182# a_2475_15206# a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3811 a_20434_14540# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3812 a_29982_12170# a_2275_12194# a_30074_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3813 VSS row_n[8] a_15318_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3814 a_20034_10162# a_2475_10186# a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3815 a_21342_3174# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3816 VDD rowon_n[1] a_11910_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3817 a_8290_13214# rowon_n[11] a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3818 a_5886_11166# a_2275_11190# a_5978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3819 a_15926_11166# a_2275_11190# a_16018_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3820 VSS row_n[8] a_5278_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3821 a_20338_7190# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3822 VSS row_n[5] a_30378_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3823 VSS row_n[1] a_31382_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3824 a_24450_13536# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3825 a_20946_10162# row_n[8] a_21438_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3826 a_2475_8178# a_1957_8178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X3827 a_5978_8154# a_2475_8178# a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3828 a_35002_3134# a_2275_3158# a_35094_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3829 a_11302_9198# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3830 a_27062_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3831 a_16322_7190# rowon_n[5] a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3832 vcm a_2275_7174# a_24050_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3833 a_22954_6146# row_n[4] a_23446_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3834 a_17326_3174# rowon_n[1] a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3835 VDD rowon_n[10] a_13918_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3836 a_33486_6508# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3837 VDD rowon_n[2] a_27974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3838 VDD rowon_n[10] a_3878_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3839 VDD rowon_n[5] a_5886_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3840 a_8898_18194# a_2275_18218# a_8990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3841 a_18938_18194# a_2275_18218# a_19030_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3842 VDD rowon_n[9] a_7894_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3843 a_20946_1126# VDD a_21438_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3844 a_26058_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3845 a_13310_15222# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3846 a_31478_1488# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3847 VDD rowon_n[0] a_3878_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3848 a_12002_17190# a_2475_17214# a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3849 a_34090_17190# a_2475_17214# a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3850 a_3270_15222# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3851 VDD VSS a_16930_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3852 a_26362_1166# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3853 a_10906_9158# row_n[7] a_11398_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3854 a_11910_5142# row_n[3] a_12402_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3855 a_4274_4178# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3856 VSS row_n[3] a_35398_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3857 a_25358_5182# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3858 a_35002_17190# row_n[15] a_35494_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3859 vcm a_2275_13198# a_35094_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3860 a_3270_8194# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3861 a_9294_2170# rowon_n[0] a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3862 a_12402_17552# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3863 a_19334_17230# rowon_n[15] a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3864 vcm a_2275_5166# a_29070_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3865 a_20338_12210# rowon_n[10] a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3866 vcm a_2275_8178# a_6982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3867 a_12914_13174# row_n[11] a_13406_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3868 a_24354_11206# rowon_n[9] a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3869 a_2874_13174# row_n[11] a_3366_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3870 a_24962_3134# row_n[1] a_25454_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3871 a_5978_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3872 a_16018_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3873 a_35494_3496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3874 a_29070_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3875 a_3878_4138# row_n[2] a_4370_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3876 VDD rowon_n[13] a_18938_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3877 VDD rowon_n[8] a_19942_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3878 a_15926_7150# row_n[5] a_16418_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3879 a_14010_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3880 a_9994_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3881 a_8290_6186# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3882 vcm a_2275_18218# a_9994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3883 a_9902_6146# a_2275_6170# a_9994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3884 a_13918_2130# row_n[0] a_14410_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3885 VSS row_n[14] a_22346_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3886 VSS row_n[13] a_35398_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3887 a_32386_12210# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3888 a_31382_9198# rowon_n[7] a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3889 a_19334_2170# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3890 vcm a_2275_3158# a_33086_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3891 a_12306_15222# rowon_n[13] a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3892 a_25054_9158# a_2475_9182# a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3893 a_30378_2170# rowon_n[0] a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3894 VSS row_n[0] a_20338_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3895 VDD VDD a_20946_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3896 VDD rowon_n[15] a_33998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3897 a_6282_14218# rowon_n[12] a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3898 a_16322_14218# rowon_n[12] a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3899 a_31478_14540# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3900 vcm a_2275_12194# a_27062_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3901 VSS row_n[9] a_3270_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3902 VSS row_n[9] a_13310_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3903 a_31078_10162# a_2475_10186# a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3904 VSS row_n[6] a_10298_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3905 a_34090_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3906 a_2874_1126# a_2275_1150# a_2966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3907 VSS row_n[2] a_11302_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3908 a_35494_13536# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3909 a_31990_10162# row_n[8] a_32482_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3910 a_14922_4138# a_2275_4162# a_15014_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3911 a_22442_5504# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3912 a_7894_13174# a_2275_13198# a_7986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3913 a_17934_13174# a_2275_13198# a_18026_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3914 VDD rowon_n[7] a_30986_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3915 VDD rowon_n[3] a_31990_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3916 VDD rowon_n[11] a_11910_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3917 a_11302_16226# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3918 a_11398_4500# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3919 a_32082_18194# a_2475_18218# a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3920 VSS row_n[1] a_3270_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3921 a_32994_18194# VDD a_33486_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3922 vcm a_2275_14202# a_33086_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3923 a_18330_12210# rowon_n[10] a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3924 VSS row_n[4] a_15318_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3925 a_10394_18556# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3926 vcm a_2275_15206# a_19030_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3927 a_5374_6508# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3928 a_5978_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3929 a_12002_4138# a_2475_4162# a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3930 vcm a_2275_15206# a_8990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3931 a_35398_11206# rowon_n[9] a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3932 a_18026_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3933 VDD rowon_n[0] a_33998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3934 a_3366_1488# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3935 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3936 a_24450_2492# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3937 a_23958_5142# a_2275_5166# a_24050_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3938 a_23046_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3939 VDD rowon_n[8] a_17934_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3940 VSS row_n[0] a_29374_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3941 a_34394_4178# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3942 a_27062_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3943 a_33390_8194# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3944 VSS row_n[3] a_7286_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3945 VSS VDD a_8290_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3946 a_18026_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3947 a_7986_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3948 a_3970_3134# a_2475_3158# a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3949 a_21342_4178# rowon_n[2] a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3950 a_35002_11166# a_2275_11190# a_35094_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3951 VSS row_n[8] a_34394_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3952 a_9390_8516# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3953 a_11302_10202# rowon_n[8] a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3954 a_9994_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3955 a_32082_2130# a_2475_2154# a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3956 a_29374_18234# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3957 VSS row_n[14] a_33390_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3958 a_27974_7150# a_2275_7174# a_28066_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3959 a_28978_3134# a_2275_3158# a_29070_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3960 a_10298_16226# rowon_n[14] a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3961 a_29470_14540# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3962 VDD rowon_n[10] a_32994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3963 a_29070_10162# a_2475_10186# a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3964 a_6890_6146# a_2275_6170# a_6982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3965 a_7382_3496# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3966 a_33998_4138# row_n[2] a_34490_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3967 vcm a_2275_4162# a_13006_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3968 a_18938_9158# a_2275_9182# a_19030_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3969 a_28066_16186# a_2475_16210# a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3970 a_20034_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3971 a_10298_3174# rowon_n[1] a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3972 VDD VDD a_31990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3973 VDD rowon_n[2] a_20946_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3974 a_28978_16186# row_n[14] a_29470_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3975 a_11910_15182# a_2275_15206# a_12002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3976 a_8990_1126# a_2475_1150# a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3977 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3978 a_15926_14178# a_2275_14202# a_16018_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3979 VDD rowon_n[4] a_11910_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3980 a_5886_14178# a_2275_14202# a_5978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3981 a_3270_9198# rowon_n[7] a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3982 a_19030_6146# a_2475_6170# a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3983 a_10298_11206# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3984 vcm a_2275_3158# a_4974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3985 VDD VSS a_9902_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3986 a_16018_9158# a_2475_9182# a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3987 a_14314_5182# rowon_n[3] a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3988 a_15318_1166# VSS a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3989 a_32994_1126# a_2275_1150# a_33086_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3990 vcm a_2275_5166# a_22042_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3991 vcm a_2275_10186# a_18026_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3992 a_19942_8154# row_n[6] a_20434_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3993 a_7894_14178# row_n[12] a_8386_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3994 a_17934_14178# row_n[12] a_18426_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3995 a_29374_12210# rowon_n[10] a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3996 vcm a_2275_10186# a_7986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3997 a_26970_10162# a_2275_10186# a_27062_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3998 VDD rowon_n[7] a_2874_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3999 a_30474_8516# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4000 VDD rowon_n[3] a_3878_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4001 VDD rowon_n[6] a_15926_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4002 vcm a_2275_16210# a_6982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4003 vcm a_2275_16210# a_17022_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4004 a_23350_3174# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4005 VDD rowon_n[1] a_13918_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4006 a_21038_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4007 VDD rowon_n[8] a_28978_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4008 a_25358_9198# rowon_n[7] a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4009 a_7986_8154# a_2475_8178# a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4010 VSS row_n[5] a_32386_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4011 VSS row_n[1] a_33390_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4012 a_13310_9198# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4013 vcm a_2275_3158# a_27062_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4014 VSS a_2161_17214# a_2275_17214# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X4015 VSS row_n[15] a_27366_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4016 a_31382_15222# rowon_n[13] a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4017 a_29070_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4018 vcm a_2275_7174# a_26058_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4019 a_24962_6146# row_n[4] a_25454_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4020 a_5978_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4021 a_16018_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4022 VDD rowon_n[5] a_7894_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4023 a_35494_6508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4024 a_28370_13214# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4025 VSS row_n[9] a_32386_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4026 vcm a_2275_9182# a_17022_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4027 a_12306_2170# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4028 a_19942_15182# a_2275_15206# a_20034_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4029 a_22954_1126# VDD a_23446_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4030 a_33486_1488# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4031 a_28066_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4032 a_14010_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4033 VSS row_n[10] a_18330_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4034 a_23046_12170# a_2475_12194# a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4035 a_31990_8154# a_2275_8178# a_32082_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4036 VDD rowon_n[0] a_5886_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4037 a_3970_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4038 VSS row_n[10] a_8290_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4039 VDD rowon_n[7] a_24962_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4040 a_28370_1166# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4041 a_27462_15544# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4042 VDD rowon_n[11] a_30986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4043 a_23958_12170# row_n[10] a_24450_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4044 a_27062_11166# a_2475_11190# a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4045 a_12914_9158# row_n[7] a_13406_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4046 a_5278_8194# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4047 a_13918_5142# row_n[3] a_14410_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4048 a_6282_4178# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4049 a_7986_10162# a_2475_10186# a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4050 a_18026_10162# a_2475_10186# a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4051 VDD rowon_n[12] a_16930_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4052 a_27974_11166# row_n[9] a_28466_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4053 VDD rowon_n[12] a_6890_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4054 vcm a_2275_8178# a_8990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4055 a_30378_16226# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4056 a_8386_10524# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4057 a_18426_10524# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4058 vcm a_2275_1150# a_31078_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4059 VDD a_2161_18218# a_2275_18218# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X4060 vcm a_2275_17214# a_21038_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4061 vcm a_2275_5166# a_30074_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4062 a_6282_17230# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4063 a_16322_17230# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4064 a_3970_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4065 vcm a_2275_16210# a_25054_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4066 a_5886_4138# row_n[2] a_6378_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4067 a_17934_7150# row_n[5] a_18426_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4068 a_8990_18194# a_2475_18218# a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4069 vcm a_2275_12194# a_12002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4070 a_15926_2130# row_n[0] a_16418_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4071 a_15926_15182# row_n[13] a_16418_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4072 a_27366_13214# rowon_n[11] a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4073 vcm a_2275_11190# a_16018_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4074 a_9390_18556# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4075 a_5886_15182# row_n[13] a_6378_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4076 vcm a_2275_11190# a_5978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4077 a_10998_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4078 a_33390_9198# rowon_n[7] a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4079 a_27366_8194# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4080 a_27062_9158# a_2475_9182# a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4081 vcm a_2275_3158# a_35094_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4082 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4083 a_19030_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4084 VSS row_n[0] a_22346_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4085 a_28978_12170# a_2275_12194# a_29070_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4086 a_32386_2170# rowon_n[0] a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4087 a_4882_1126# a_2275_1150# a_4974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4088 a_19030_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4089 VSS row_n[2] a_13310_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4090 VDD rowon_n[9] a_26970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4091 VSS row_n[6] a_12306_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4092 a_26058_2130# a_2475_2154# a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4093 a_24450_5504# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4094 VDD rowon_n[7] a_32994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4095 VDD rowon_n[3] a_33998_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4096 VSS VDD a_25358_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4097 a_22346_15222# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4098 a_2966_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4099 a_26362_14218# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4100 a_2161_10186# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4101 a_20946_7150# a_2275_7174# a_21038_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4102 VSS a_2161_5166# a_2275_5166# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X4103 a_21950_3134# a_2275_3158# a_22042_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4104 a_15318_17230# rowon_n[15] a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4105 a_31078_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4106 a_34090_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4107 a_5278_17230# rowon_n[15] a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4108 a_30986_15182# a_2275_15206# a_31078_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4109 a_11910_9158# a_2275_9182# a_12002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4110 a_12002_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4111 a_21438_17552# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4112 a_9294_16226# rowon_n[14] a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4113 VSS row_n[11] a_6282_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4114 VSS row_n[11] a_16322_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4115 a_21038_13174# a_2475_13198# a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4116 a_19334_6186# rowon_n[4] a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4117 a_31382_6186# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4118 VSS row_n[1] a_5278_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4119 a_13406_4500# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4120 a_25454_16548# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4121 a_35002_14178# a_2275_14202# a_35094_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4122 a_21950_13174# row_n[11] a_22442_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4123 VSS row_n[5] a_4274_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4124 a_16018_11166# a_2475_11190# a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4125 VSS row_n[4] a_17326_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4126 a_5978_11166# a_2475_11190# a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4127 a_7382_6508# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4128 VDD rowon_n[13] a_4882_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4129 VDD rowon_n[13] a_14922_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4130 a_7986_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4131 a_14010_4138# a_2475_4162# a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4132 a_5278_12210# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4133 a_15318_12210# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4134 vcm a_2275_12194# a_20034_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4135 a_16418_11528# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4136 a_26970_1126# a_2275_1150# a_27062_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4137 a_25966_5142# a_2275_5166# a_26058_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4138 a_6378_11528# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4139 a_3878_8154# a_2275_8178# a_3970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4140 vcm a_2275_6170# a_9994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4141 a_5374_1488# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4142 a_14314_18234# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4143 a_4274_18234# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4144 vcm a_2275_17214# a_32082_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4145 a_35398_8194# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4146 a_4370_14540# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4147 a_14410_14540# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4148 VSS row_n[3] a_9294_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4149 a_14922_10162# row_n[8] a_15414_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4150 a_23046_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4151 a_4882_10162# row_n[8] a_5374_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4152 a_23350_4178# rowon_n[2] a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4153 a_2161_8178# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X4154 VSS row_n[5] a_26362_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4155 a_3878_16186# row_n[14] a_4370_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4156 a_13918_16186# row_n[14] a_14410_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4157 a_25358_14218# rowon_n[12] a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4158 a_1957_13198# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4159 a_34090_2130# a_2475_2154# a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4160 vcm a_2275_1150# a_2966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4161 a_8898_6146# a_2275_6170# a_8990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4162 a_9390_3496# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4163 vcm a_2275_4162# a_15014_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4164 a_26058_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4165 a_23350_17230# rowon_n[15] a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4166 a_26970_13174# a_2275_13198# a_27062_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4167 a_29982_3134# a_2275_3158# a_30074_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4168 a_22042_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4169 a_11302_7190# rowon_n[5] a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4170 a_12306_3174# rowon_n[1] a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4171 VSS row_n[11] a_24354_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4172 a_21342_10202# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4173 VDD rowon_n[2] a_22954_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4174 a_14314_12210# rowon_n[10] a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4175 VDD rowon_n[4] a_13918_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4176 a_21038_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4177 a_4274_12210# rowon_n[10] a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4178 a_11910_10162# a_2275_10186# a_12002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4179 a_19430_17552# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4180 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4181 VDD rowon_n[13] a_22954_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4182 a_19030_13174# a_2475_13198# a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4183 a_20434_12532# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4184 VDD VSS a_11910_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4185 a_21342_1166# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4186 a_8290_11206# rowon_n[9] a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4187 VSS VDD a_31382_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4188 VSS row_n[3] a_30378_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4189 a_20338_5182# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4190 a_24450_11528# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4191 a_5978_6146# a_2475_6170# a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4192 a_35002_1126# a_2275_1150# a_35094_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4193 a_4274_2170# rowon_n[0] a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4194 a_18026_9158# a_2475_9182# a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4195 a_16322_5182# rowon_n[3] a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4196 a_17326_1166# VSS a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4197 vcm a_2275_5166# a_24050_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4198 a_35398_17230# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4199 VDD rowon_n[8] a_13918_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4200 a_32482_8516# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4201 VDD rowon_n[8] a_3878_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4202 VDD rowon_n[3] a_5886_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4203 VSS row_n[15] a_12306_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4204 a_8898_16186# a_2275_16210# a_8990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4205 a_18938_16186# a_2275_16210# a_19030_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4206 a_19942_3134# row_n[1] a_20434_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4207 a_13310_13214# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4208 a_30474_3496# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4209 a_12002_15182# a_2475_15206# a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4210 a_34090_15182# a_2475_15206# a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4211 a_3270_13214# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4212 vcm a_2275_12194# a_31078_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4213 a_25358_3174# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4214 a_10906_7150# row_n[5] a_11398_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4215 VSS row_n[1] a_35398_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4216 VDD rowon_n[1] a_15926_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4217 a_35002_15182# row_n[13] a_35494_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4218 vcm a_2275_11190# a_35094_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4219 a_27366_9198# rowon_n[7] a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4220 a_9994_8154# a_2475_8178# a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4221 VSS row_n[5] a_34394_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4222 a_3270_6186# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4223 a_12402_15544# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4224 a_19334_15222# rowon_n[13] a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4225 a_20338_10202# rowon_n[8] a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4226 a_15318_9198# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4227 vcm a_2275_7174# a_28066_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4228 vcm a_2275_3158# a_29070_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4229 a_21038_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4230 vcm a_2275_6170# a_6982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4231 a_12914_11166# row_n[9] a_13406_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4232 vcm a_2275_9182# a_19030_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4233 VSS a_2161_12194# a_2275_12194# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X4234 a_2874_11166# row_n[9] a_3366_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4235 a_24962_1126# VDD a_25454_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4236 a_14314_2170# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4237 a_25054_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4238 a_20034_9158# a_2475_9182# a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4239 a_33998_8154# a_2275_8178# a_34090_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4240 a_35494_1488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4241 VDD rowon_n[0] a_7894_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4242 VDD rowon_n[11] a_18938_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4243 a_19942_10162# a_2275_10186# a_20034_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4244 a_14922_9158# row_n[7] a_15414_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4245 VDD rowon_n[7] a_26970_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4246 a_15926_5142# row_n[3] a_16418_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4247 a_8290_4178# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4248 a_21342_18234# VDD a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4249 vcm a_2275_16210# a_9994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4250 a_9902_4138# a_2275_4162# a_9994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4251 a_34394_17230# rowon_n[15] a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4252 VSS row_n[12] a_22346_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4253 VSS row_n[11] a_35398_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4254 a_32386_10202# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4255 a_22954_17190# a_2275_17214# a_23046_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4256 vcm a_2275_1150# a_33086_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4257 a_12306_13214# rowon_n[11] a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4258 a_7894_4138# row_n[2] a_8386_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4259 VDD rowon_n[14] a_20946_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4260 VDD rowon_n[13] a_33998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4261 a_26970_14178# row_n[12] a_27462_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4262 a_31478_12532# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4263 vcm a_2275_10186# a_27062_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4264 a_13918_12170# a_2275_12194# a_14010_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4265 VSS row_n[4] a_10298_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4266 a_3878_12170# a_2275_12194# a_3970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4267 a_35494_11528# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4268 VDD rowon_n[5] a_30986_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4269 a_17934_2130# row_n[0] a_18426_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4270 a_33390_18234# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4271 VDD rowon_n[9] a_11910_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4272 a_29374_8194# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4273 VSS VDD a_10298_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4274 a_13006_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4275 a_29070_9158# a_2475_9182# a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4276 vcm a_2275_18218# a_28066_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4277 a_32082_16186# a_2475_16210# a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4278 a_11302_14218# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4279 VSS row_n[0] a_24354_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4280 a_18330_10202# rowon_n[8] a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4281 a_34394_2170# rowon_n[0] a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4282 VSS VDD a_3270_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4283 a_32994_16186# row_n[14] a_33486_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4284 a_19030_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4285 VSS row_n[6] a_14314_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4286 a_28066_2130# a_2475_2154# a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4287 VSS row_n[2] a_15318_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4288 vcm a_2275_8178# a_32082_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4289 a_18938_17190# row_n[15] a_19430_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4290 a_10394_16548# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4291 vcm a_2275_13198# a_19030_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4292 a_4370_8516# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4293 a_5978_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4294 a_8898_17190# row_n[15] a_9390_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4295 vcm a_2275_13198# a_8990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4296 a_4974_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4297 a_23958_3134# a_2275_3158# a_24050_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4298 VDD a_2161_9182# a_2275_9182# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X4299 a_22954_7150# a_2275_7174# a_23046_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4300 a_23046_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4301 a_33086_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4302 a_13918_9158# a_2275_9182# a_14010_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4303 a_33390_6186# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4304 VSS row_n[1] a_7286_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4305 a_15414_4500# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4306 a_33390_12210# rowon_n[10] a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4307 a_30986_10162# a_2275_10186# a_31078_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4308 a_3970_1126# a_2475_1150# a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4309 a_32386_18234# VDD a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4310 a_9390_6508# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4311 a_9994_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4312 a_28978_1126# a_2275_1150# a_29070_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4313 a_29374_16226# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4314 VSS row_n[12] a_33390_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4315 a_27974_5142# a_2275_5166# a_28066_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4316 a_20946_18194# a_2275_18218# a_21038_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4317 a_33998_17190# a_2275_17214# a_34090_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4318 a_10298_14218# rowon_n[12] a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4319 a_29470_12532# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4320 VDD rowon_n[8] a_32994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4321 a_5886_8154# a_2275_8178# a_5978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4322 a_7382_1488# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4323 a_6890_4138# a_2275_4162# a_6982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4324 a_26458_8516# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4325 a_28066_14178# a_2475_14202# a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4326 a_10998_9158# a_2475_9182# a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4327 a_10298_1166# VSS a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4328 a_28466_18556# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4329 VDD rowon_n[14] a_31990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4330 a_11910_13174# a_2275_13198# a_12002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4331 VDD rowon_n[6] a_10906_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4332 VSS row_n[5] a_28370_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4333 a_19030_4138# a_2475_4162# a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4334 a_1957_7174# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4335 vcm a_2275_1150# a_4974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4336 a_20338_9198# rowon_n[7] a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4337 a_2966_8154# a_2475_8178# a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4338 a_13310_7190# rowon_n[5] a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4339 vcm a_2275_3158# a_22042_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4340 a_14314_3174# rowon_n[1] a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4341 a_24050_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4342 vcm a_2275_7174# a_21038_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4343 a_31078_7150# a_2475_7174# a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4344 a_19942_6146# row_n[4] a_20434_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4345 a_7894_12170# row_n[10] a_8386_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4346 a_17934_12170# row_n[10] a_18426_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4347 a_29374_10202# rowon_n[8] a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4348 VDD rowon_n[5] a_2874_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4349 a_30474_6508# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4350 vcm a_2275_9182# a_12002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4351 VDD rowon_n[4] a_15926_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4352 a_16930_18194# VDD a_17422_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4353 vcm a_2275_14202# a_6982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4354 vcm a_2275_14202# a_17022_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4355 a_23046_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4356 a_6890_18194# VDD a_7382_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4357 VDD rowon_n[7] a_19942_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4358 VDD VSS a_13918_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4359 a_23350_1166# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4360 vcm a_2275_17214# a_15014_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4361 a_21038_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4362 a_7986_6146# a_2475_6170# a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4363 VSS VDD a_33390_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4364 a_6282_2170# rowon_n[0] a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4365 VSS row_n[3] a_32386_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4366 vcm a_2275_17214# a_4974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4367 vcm a_2275_1150# a_27062_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4368 VSS a_2161_15206# a_2275_15206# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X4369 VSS row_n[13] a_27366_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4370 a_31382_13214# rowon_n[11] a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4371 a_24354_12210# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4372 vcm a_2275_5166# a_26058_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4373 vcm a_2275_8178# a_3970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4374 a_34490_8516# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4375 VDD rowon_n[3] a_7894_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4376 a_28370_11206# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4377 a_19942_13174# a_2275_13198# a_20034_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4378 VDD rowon_n[15] a_25966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4379 a_14010_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4380 a_23446_14540# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4381 a_32994_12170# a_2275_12194# a_33086_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4382 VSS row_n[8] a_18330_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4383 a_23046_10162# a_2475_10186# a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4384 a_31990_6146# a_2275_6170# a_32082_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4385 a_32482_3496# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4386 a_3970_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4387 a_8898_11166# a_2275_11190# a_8990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4388 a_18938_11166# a_2275_11190# a_19030_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4389 VSS row_n[8] a_8290_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4390 VDD rowon_n[5] a_24962_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4391 a_31990_18194# a_2275_18218# a_32082_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4392 a_27462_13536# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4393 VDD rowon_n[9] a_30986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4394 a_23958_10162# row_n[8] a_24450_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4395 VSS row_n[7] a_19334_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4396 a_12914_7150# row_n[5] a_13406_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4397 a_5278_6186# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4398 a_29374_9198# rowon_n[7] a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4399 VDD rowon_n[10] a_16930_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4400 a_10906_2130# row_n[0] a_11398_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4401 VDD rowon_n[10] a_6890_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4402 vcm a_2275_6170# a_8990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4403 a_30378_14218# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4404 a_22346_8194# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4405 a_24050_18194# a_2475_18218# a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4406 VDD a_2161_16210# a_2275_16210# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X4407 a_16322_15222# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4408 vcm a_2275_15206# a_21038_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4409 a_22042_9158# a_2475_9182# a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4410 a_16322_2170# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4411 vcm a_2275_3158# a_30074_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4412 VSS VDD a_9294_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4413 a_15014_17190# a_2475_17214# a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4414 a_6282_15222# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4415 a_19430_9520# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4416 a_24962_18194# VDD a_25454_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4417 a_4974_17190# a_2475_17214# a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4418 vcm a_2275_14202# a_25054_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4419 VDD rowon_n[7] a_28978_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4420 a_17934_5142# row_n[3] a_18426_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4421 a_15414_17552# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4422 a_8990_16186# a_2475_16210# a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4423 vcm a_2275_10186# a_12002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4424 a_21038_2130# a_2475_2154# a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4425 a_5374_17552# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4426 a_11910_14178# row_n[12] a_12402_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4427 a_15926_13174# row_n[11] a_16418_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4428 a_27366_11206# rowon_n[9] a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4429 a_9390_16548# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4430 a_5886_13174# row_n[11] a_6378_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4431 a_27366_6186# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4432 vcm a_2275_1150# a_35094_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4433 a_19030_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4434 vcm a_2275_18218# a_2966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4435 vcm a_2275_18218# a_13006_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4436 VSS row_n[15] a_21342_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4437 VSS row_n[4] a_12306_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4438 VDD rowon_n[5] a_32994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4439 VSS row_n[14] a_25358_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4440 a_22346_13214# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4441 a_2966_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4442 a_15014_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4443 a_21950_1126# a_2275_1150# a_22042_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4444 VSS a_2161_3158# a_2275_3158# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X4445 a_20946_5142# a_2275_5166# a_21038_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4446 a_30074_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4447 a_15318_15222# rowon_n[13] a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4448 VDD rowon_n[0] a_30986_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4449 a_31078_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4450 a_34090_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4451 a_5278_15222# rowon_n[13] a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4452 a_30986_13174# a_2275_13198# a_31078_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4453 VDD VDD a_23958_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4454 a_12002_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4455 a_21438_15544# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4456 a_9294_14218# rowon_n[12] a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4457 VSS row_n[9] a_6282_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4458 VSS row_n[9] a_16322_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4459 a_21038_11166# a_2475_11190# a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4460 a_18330_8194# rowon_n[6] a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4461 a_30378_8194# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4462 VSS VDD a_5278_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4463 a_31382_4178# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4464 a_19334_4178# rowon_n[2] a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4465 a_21950_11166# row_n[9] a_22442_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4466 VSS row_n[3] a_4274_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4467 VSS row_n[2] a_17326_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4468 vcm a_2275_8178# a_34090_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4469 VDD rowon_n[11] a_4882_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4470 VDD rowon_n[11] a_14922_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4471 a_6982_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4472 VSS row_n[5] a_21342_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4473 a_7986_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4474 a_19942_14178# row_n[12] a_20434_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4475 a_5278_10202# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4476 a_15318_10202# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4477 vcm a_2275_10186# a_20034_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4478 a_24962_7150# a_2275_7174# a_25054_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4479 a_25966_3134# a_2275_3158# a_26058_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4480 a_3970_12170# a_2475_12194# a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4481 a_14010_12170# a_2475_12194# a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4482 a_35094_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4483 a_3878_6146# a_2275_6170# a_3970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4484 a_4370_3496# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4485 VDD rowon_n[2] a_18938_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4486 vcm a_2275_4162# a_9994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4487 a_14314_16226# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4488 a_15926_9158# a_2275_9182# a_16018_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4489 a_30986_4138# row_n[2] a_31478_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4490 a_13006_18194# a_2475_18218# a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4491 a_35094_18194# a_2475_18218# a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4492 a_4274_16226# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4493 vcm a_2275_15206# a_32082_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4494 a_35398_6186# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4495 VSS row_n[1] a_9294_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4496 a_17422_4500# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4497 a_2966_18194# a_2475_18218# a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4498 a_4370_12532# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4499 a_14410_12532# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4500 a_13406_18556# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4501 a_3366_18556# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4502 VSS row_n[3] a_26362_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4503 a_1957_11190# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4504 a_1957_1150# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X4505 a_26058_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4506 a_7894_8154# a_2275_8178# a_7986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4507 a_9390_1488# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4508 a_8898_4138# a_2275_4162# a_8990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4509 a_28466_8516# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4510 VSS row_n[15] a_19334_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4511 a_23350_15222# rowon_n[13] a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4512 VSS row_n[10] a_20338_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4513 a_29982_1126# a_2275_1150# a_30074_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4514 a_13006_9158# a_2475_9182# a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4515 a_11302_5182# rowon_n[3] a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4516 a_12306_1166# VSS a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4517 VSS row_n[9] a_24354_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4518 a_26458_3496# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4519 a_14314_10202# rowon_n[8] a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4520 VDD rowon_n[6] a_12914_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4521 a_4274_10202# rowon_n[8] a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4522 a_19430_15544# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4523 VDD rowon_n[11] a_22954_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4524 a_19030_11166# a_2475_11190# a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4525 a_20434_10524# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4526 a_20338_3174# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4527 VSS row_n[1] a_30378_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4528 VDD rowon_n[1] a_10906_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4529 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4530 a_22346_9198# rowon_n[7] a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4531 a_4974_8154# a_2475_8178# a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4532 a_5978_4138# a_2475_4162# a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4533 VDD VDD a_35002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4534 a_10298_9198# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4535 vcm a_2275_7174# a_23046_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4536 vcm a_2275_3158# a_24050_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4537 a_16322_3174# rowon_n[1] a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4538 a_35398_15222# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4539 a_33086_7150# a_2475_7174# a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4540 a_32482_6508# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4541 vcm a_2275_9182# a_14010_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4542 VSS row_n[13] a_12306_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4543 a_8898_14178# a_2275_14202# a_8990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4544 a_18938_14178# a_2275_14202# a_19030_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4545 a_19942_1126# en_bit_n[0] a_20434_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4546 a_25054_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4547 a_13310_11206# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4548 a_30474_1488# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4549 a_34490_17552# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4550 a_30986_14178# row_n[12] a_31478_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4551 a_12002_13174# a_2475_13198# a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4552 a_34090_13174# a_2475_13198# a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4553 a_3270_11206# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4554 vcm a_2275_10186# a_31078_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4555 VDD VSS a_15926_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4556 a_25358_1166# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4557 VDD rowon_n[0] a_2874_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4558 a_9902_9158# row_n[7] a_10394_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4559 VDD rowon_n[7] a_21950_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4560 a_10906_5142# row_n[3] a_11398_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4561 VDD rowon_n[15] a_10906_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4562 a_35002_13174# row_n[11] a_35494_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4563 a_9994_6146# a_2475_6170# a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4564 a_8290_2170# rowon_n[0] a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4565 a_3270_4178# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4566 VSS row_n[3] a_34394_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4567 a_12402_13536# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4568 a_19334_13214# rowon_n[11] a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4569 vcm a_2275_1150# a_29070_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4570 vcm a_2275_5166# a_28066_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4571 vcm a_2275_8178# a_5978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4572 vcm a_2275_4162# a_6982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4573 a_2475_7174# a_1957_7174# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X4574 VSS a_2161_10186# a_2275_10186# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X4575 a_33998_6146# a_2275_6170# a_34090_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4576 a_34490_3496# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4577 a_2874_4138# row_n[2] a_3366_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4578 VDD rowon_n[9] a_18938_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4579 a_14922_7150# row_n[5] a_15414_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4580 VDD rowon_n[5] a_26970_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4581 a_2475_18218# a_1957_18218# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X4582 a_14010_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4583 a_9902_18194# VDD a_10394_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4584 a_21342_16226# rowon_n[14] a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4585 a_34394_15222# rowon_n[13] a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4586 vcm a_2275_14202# a_9994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4587 VSS row_n[10] a_31382_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4588 a_3970_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4589 VDD rowon_n[0] a_24962_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4590 a_12914_2130# row_n[0] a_13406_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4591 VSS row_n[9] a_35398_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4592 a_24354_8194# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4593 a_22954_15182# a_2275_15206# a_23046_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4594 a_18330_2170# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4595 a_17022_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4596 VDD rowon_n[12] a_29982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4597 a_26058_12170# a_2475_12194# a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4598 a_12306_11206# rowon_n[9] a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4599 a_24050_9158# a_2475_9182# a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4600 a_6982_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4601 VDD rowon_n[11] a_33998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4602 a_26970_12170# row_n[10] a_27462_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4603 a_31478_10524# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4604 a_23046_2130# a_2475_2154# a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4605 VSS row_n[2] a_10298_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4606 VDD rowon_n[3] a_30986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4607 a_33390_16226# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4608 a_29374_6186# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4609 VSS row_n[14] a_10298_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4610 a_9294_17230# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4611 a_19334_17230# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4612 vcm a_2275_17214# a_24050_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4613 a_7286_9198# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4614 vcm a_2275_16210# a_28066_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4615 a_32082_14178# a_2475_14202# a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4616 a_10394_4500# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4617 a_14922_18194# a_2275_18218# a_15014_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4618 a_32482_18556# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4619 a_4882_18194# a_2275_18218# a_4974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4620 VSS row_n[4] a_14314_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4621 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4622 vcm a_2275_6170# a_32082_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4623 a_18938_15182# row_n[13] a_19430_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4624 vcm a_2275_11190# a_19030_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4625 a_4370_6508# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4626 a_8898_15182# row_n[13] a_9390_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4627 vcm a_2275_11190# a_8990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4628 a_6890_9158# row_n[7] a_7382_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4629 a_4974_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4630 a_23958_1126# a_2275_1150# a_24050_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4631 a_17022_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4632 a_33086_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4633 a_22954_5142# a_2275_5166# a_23046_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4634 VDD rowon_n[0] a_32994_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4635 a_21438_8516# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4636 VSS row_n[10] a_29374_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4637 VSS VDD a_7286_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4638 a_16018_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4639 a_33390_4178# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4640 a_34090_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4641 a_33390_10202# rowon_n[8] a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4642 a_12002_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4643 VSS VDD a_28370_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4644 a_32386_16226# rowon_n[14] a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4645 VDD rowon_n[12] a_27974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4646 a_8990_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4647 VSS row_n[5] a_23350_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4648 a_9994_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4649 a_29374_14218# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4650 a_27974_3134# a_2275_3158# a_28066_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4651 a_20946_16186# a_2275_16210# a_21038_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4652 a_33998_15182# a_2275_15206# a_34090_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4653 a_29470_10524# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4654 a_5886_6146# a_2275_6170# a_5978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4655 a_32994_4138# row_n[2] a_33486_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4656 a_4974_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4657 a_15014_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4658 a_17934_9158# a_2275_9182# a_18026_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4659 a_26458_6508# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4660 a_28466_16548# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4661 a_16930_2130# a_2275_2154# a_17022_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4662 VDD rowon_n[4] a_10906_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4663 a_8290_12210# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4664 a_18330_12210# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4665 vcm a_2275_12194# a_23046_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4666 VSS row_n[3] a_28370_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4667 VSS row_n[6] a_6282_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4668 a_1957_5166# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4669 a_17326_18234# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4670 vcm a_2275_18218# a_22042_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4671 a_7286_18234# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4672 a_2966_6146# a_2475_6170# a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4673 a_7382_14540# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4674 a_17422_14540# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4675 a_13310_5182# rowon_n[3] a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4676 a_14314_1166# VSS a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4677 vcm a_2275_1150# a_22042_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4678 a_26058_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4679 a_15014_9158# a_2475_9182# a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4680 a_28466_3496# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4681 a_31078_5142# a_2475_5166# a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4682 vcm a_2275_5166# a_21038_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4683 a_7894_10162# row_n[8] a_8386_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4684 a_17934_10162# row_n[8] a_18426_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4685 VDD rowon_n[3] a_2874_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4686 a_16930_16186# row_n[14] a_17422_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4687 a_6890_16186# row_n[14] a_7382_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4688 VDD rowon_n[5] a_19942_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4689 VDD rowon_n[1] a_12914_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4690 a_26362_17230# rowon_n[15] a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4691 vcm a_2275_15206# a_15014_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4692 VSS row_n[1] a_32386_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4693 a_7986_4138# a_2475_4162# a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4694 vcm a_2275_15206# a_4974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4695 a_24354_9198# rowon_n[7] a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4696 a_6982_8154# a_2475_8178# a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4697 VSS row_n[11] a_27366_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4698 a_31382_11206# rowon_n[9] a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4699 a_24354_10202# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4700 vcm a_2275_7174# a_25054_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4701 vcm a_2275_3158# a_26058_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4702 a_35094_7150# a_2475_7174# a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4703 vcm a_2275_6170# a_3970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4704 a_34490_6508# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4705 a_17326_12210# rowon_n[10] a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4706 vcm a_2275_9182# a_16018_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4707 a_2475_1150# a_1957_1150# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X4708 a_7286_12210# rowon_n[10] a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4709 a_27062_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4710 a_11302_2170# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4711 VDD rowon_n[13] a_25966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4712 a_14010_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4713 a_23446_12532# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4714 a_30986_8154# a_2275_8178# a_31078_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4715 a_32482_1488# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4716 a_31990_4138# a_2275_4162# a_32082_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4717 a_3970_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4718 VDD rowon_n[7] a_23958_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4719 VDD rowon_n[3] a_24962_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4720 a_31990_16186# a_2275_16210# a_32082_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4721 a_27462_11528# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4722 a_12914_5142# row_n[3] a_13406_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4723 a_5278_4178# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4724 a_25358_18234# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4725 VDD rowon_n[8] a_16930_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4726 VDD rowon_n[8] a_6890_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4727 vcm a_2275_8178# a_7986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4728 vcm a_2275_4162# a_8990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4729 VSS row_n[15] a_5278_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4730 VSS row_n[15] a_15318_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4731 a_20034_17190# a_2475_17214# a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4732 a_22346_6186# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4733 a_24050_16186# a_2475_16210# a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4734 VDD a_2161_14202# a_2275_14202# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X4735 a_16322_13214# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4736 vcm a_2275_13198# a_21038_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4737 a_5278_7190# rowon_n[5] a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4738 vcm a_2275_1150# a_30074_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4739 a_20946_17190# row_n[15] a_21438_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4740 VSS row_n[14] a_9294_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4741 a_15014_15182# a_2475_15206# a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4742 a_6282_13214# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4743 vcm a_2275_12194# a_34090_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4744 a_19430_7512# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4745 a_24962_16186# row_n[14] a_25454_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4746 a_4974_15182# a_2475_15206# a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4747 VDD rowon_n[5] a_28978_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4748 a_4882_4138# row_n[2] a_5374_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4749 a_15414_15544# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4750 a_8990_14178# a_2475_14202# a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4751 a_11910_12170# row_n[10] a_12402_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4752 VDD VDD a_7894_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4753 a_5374_15544# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4754 VDD rowon_n[0] a_26970_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4755 a_2475_13198# a_1957_13198# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X4756 a_15926_11166# row_n[9] a_16418_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4757 a_14922_2130# row_n[0] a_15414_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4758 a_5886_11166# row_n[9] a_6378_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4759 a_26362_8194# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4760 a_27366_4178# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4761 a_28066_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4762 a_22954_10162# a_2275_10186# a_23046_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4763 a_31382_2170# rowon_n[0] a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4764 VSS row_n[2] a_12306_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4765 a_24354_18234# VDD a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4766 vcm a_2275_16210# a_2966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4767 vcm a_2275_16210# a_13006_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4768 VSS row_n[13] a_21342_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4769 a_25054_2130# a_2475_2154# a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4770 a_26970_4138# row_n[2] a_27462_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4771 VDD rowon_n[3] a_32994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4772 VSS row_n[12] a_25358_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4773 a_22346_11206# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4774 a_2966_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4775 a_25966_17190# a_2275_17214# a_26058_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4776 a_30074_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4777 a_19942_7150# a_2275_7174# a_20034_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4778 a_20946_3134# a_2275_3158# a_21038_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4779 VDD rowon_n[15] a_19942_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4780 a_15318_13214# rowon_n[11] a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4781 a_9294_9198# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4782 a_30074_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4783 a_31078_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4784 a_34090_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4785 a_5278_13214# rowon_n[11] a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4786 a_10906_9158# a_2275_9182# a_10998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4787 VDD rowon_n[14] a_23958_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4788 a_12002_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4789 a_21438_13536# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4790 a_18330_6186# rowon_n[4] a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4791 a_30378_6186# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4792 VSS row_n[1] a_4274_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4793 a_12402_4500# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4794 a_16930_12170# a_2275_12194# a_17022_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4795 a_6890_12170# a_2275_12194# a_6982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4796 VSS row_n[10] a_14314_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4797 vcm a_2275_6170# a_34090_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4798 VSS row_n[10] a_4274_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4799 VDD rowon_n[9] a_4882_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4800 VDD rowon_n[9] a_14922_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4801 a_6982_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4802 VSS row_n[3] a_21342_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4803 VSS VDD a_13310_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4804 a_19942_12170# row_n[10] a_20434_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4805 a_8898_9158# row_n[7] a_9390_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4806 a_25966_1126# a_2275_1150# a_26058_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4807 a_24962_5142# a_2275_5166# a_25054_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4808 VSS VDD a_3270_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4809 a_31078_17190# a_2475_17214# a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4810 a_3970_10162# a_2475_10186# a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4811 a_14010_10162# a_2475_10186# a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4812 a_2874_8154# a_2275_8178# a_2966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4813 a_4370_1488# en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4814 a_3878_4138# a_2275_4162# a_3970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4815 a_35094_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4816 VDD rowon_n[12] a_12914_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4817 a_14314_14218# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4818 a_23446_8516# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4819 a_31990_17190# row_n[15] a_32482_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4820 a_13006_16186# a_2475_16210# a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4821 a_35094_16186# a_2475_16210# a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4822 VDD rowon_n[12] a_2874_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4823 a_4274_14218# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4824 vcm a_2275_13198# a_32082_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4825 VSS VDD a_9294_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4826 a_35398_4178# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4827 a_2966_16186# a_2475_16210# a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4828 a_4370_10524# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4829 a_14410_10524# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4830 a_18026_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4831 a_21438_3496# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4832 a_13406_16548# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4833 a_3366_16548# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4834 VSS row_n[5] a_25358_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4835 VSS row_n[1] a_26362_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4836 a_35398_7190# rowon_n[5] a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4837 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4838 a_26058_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4839 VSS row_n[7] a_16322_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4840 a_7894_6146# a_2275_6170# a_7986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4841 a_28466_6508# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4842 a_35002_4138# row_n[2] a_35494_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4843 VSS row_n[13] a_19334_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4844 a_23350_13214# rowon_n[11] a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4845 VSS row_n[8] a_20338_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4846 a_20946_11166# a_2275_11190# a_21038_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4847 a_11302_3174# rowon_n[1] a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4848 a_33998_10162# a_2275_10186# a_34090_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4849 a_26458_1488# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4850 a_35398_18234# VDD a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4851 a_18938_2130# a_2275_2154# a_19030_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4852 VDD rowon_n[15] a_17934_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4853 a_24962_12170# a_2275_12194# a_25054_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4854 VDD rowon_n[4] a_12914_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4855 a_20034_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4856 a_16418_9520# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4857 VSS row_n[6] a_8290_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4858 a_23958_18194# a_2275_18218# a_24050_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4859 a_19430_13536# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4860 VDD rowon_n[9] a_22954_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4861 VDD VSS a_10906_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4862 VSS VDD a_30378_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4863 VSS row_n[15] a_34394_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4864 a_2161_7174# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4865 a_4974_6146# a_2475_6170# a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4866 a_3270_2170# rowon_n[0] a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4867 VDD rowon_n[14] a_35002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4868 a_17022_9158# a_2475_9182# a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4869 a_16322_1166# VSS a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4870 vcm a_2275_1150# a_24050_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4871 vcm a_2275_5166# a_23046_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4872 a_11302_17230# rowon_n[15] a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4873 a_35398_13214# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4874 a_33086_5142# a_2475_5166# a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4875 a_29070_17190# a_2475_17214# a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4876 VSS row_n[11] a_12306_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4877 a_30074_12170# a_2475_12194# a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4878 a_16018_2130# a_2475_2154# a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4879 a_34490_15544# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4880 a_30986_12170# row_n[10] a_31478_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4881 a_12002_11166# a_2475_11190# a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4882 a_34090_11166# a_2475_11190# a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4883 a_9902_7150# row_n[5] a_10394_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4884 VDD rowon_n[5] a_21950_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4885 VSS row_n[1] a_34394_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4886 VDD rowon_n[13] a_10906_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4887 a_35002_11166# row_n[9] a_35494_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4888 a_26362_9198# rowon_n[7] a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4889 a_8990_8154# a_2475_8178# a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4890 a_9994_4138# a_2475_4162# a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4891 a_12402_11528# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4892 a_19334_11206# rowon_n[9] a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4893 VDD rowon_n[0] a_19942_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4894 vcm a_2275_3158# a_28066_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4895 vcm a_2275_6170# a_5978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4896 a_10298_18234# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4897 vcm a_2275_9182# a_18026_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4898 a_2475_5166# a_1957_5166# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X4899 a_25358_2170# rowon_n[0] a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4900 a_13310_2170# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4901 a_32994_8154# a_2275_8178# a_33086_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4902 a_29070_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4903 a_33998_4138# a_2275_4162# a_34090_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4904 a_15318_8194# rowon_n[6] a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4905 vcm a_2275_17214# a_18026_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4906 VDD rowon_n[7] a_25966_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4907 a_14922_5142# row_n[3] a_15414_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4908 vcm a_2275_2154# a_17022_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4909 VDD rowon_n[3] a_26970_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4910 vcm a_2275_17214# a_7986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4911 VDD rowon_n[6] a_4882_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4912 a_9902_16186# row_n[14] a_10394_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4913 a_21342_14218# rowon_n[12] a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4914 a_34394_13214# rowon_n[11] a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4915 a_27366_12210# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4916 VSS row_n[8] a_31382_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4917 a_22042_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4918 a_31990_11166# a_2275_11190# a_32082_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4919 a_24354_6186# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4920 a_22954_13174# a_2275_13198# a_23046_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4921 VDD rowon_n[15] a_28978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4922 a_17022_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4923 a_26458_14540# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4924 VDD rowon_n[10] a_29982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4925 a_26058_10162# a_2475_10186# a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4926 a_7286_7190# rowon_n[5] a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4927 a_6982_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4928 VDD rowon_n[9] a_33998_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4929 a_26970_10162# row_n[8] a_27462_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4930 VSS VDD a_32386_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4931 VDD rowon_n[0] a_28978_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4932 a_19430_2492# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4933 a_33390_14218# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4934 a_29374_4178# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4935 a_27062_18194# a_2475_18218# a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4936 vcm a_2275_15206# a_24050_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4937 VSS row_n[12] a_10298_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4938 a_12002_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4939 a_28370_8194# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4940 a_18026_17190# a_2475_17214# a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4941 a_9294_15222# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4942 a_19334_15222# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4943 a_27974_18194# VDD a_28466_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4944 a_7986_17190# a_2475_17214# a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4945 a_10906_17190# a_2275_17214# a_10998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4946 vcm a_2275_14202# a_28066_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4947 a_14922_16186# a_2275_16210# a_15014_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4948 a_32482_16548# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4949 a_33390_2170# rowon_n[0] a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4950 a_10998_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4951 a_4882_16186# a_2275_16210# a_4974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4952 a_27062_2130# a_2475_2154# a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4953 VSS row_n[2] a_14314_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4954 a_8386_17552# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4955 a_18426_17552# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4956 vcm a_2275_8178# a_31078_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4957 a_17326_7190# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4958 vcm a_2275_4162# a_32082_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4959 a_18938_13174# row_n[11] a_19430_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4960 a_28978_4138# row_n[2] a_29470_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4961 a_8898_13174# row_n[11] a_9390_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4962 a_3970_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4963 a_6890_7150# row_n[5] a_7382_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4964 a_4974_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4965 a_33086_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4966 a_22954_3134# a_2275_3158# a_23046_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4967 a_2161_16210# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X4968 a_32082_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4969 a_12914_9158# a_2275_9182# a_13006_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4970 a_21438_6508# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4971 a_30074_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4972 VSS row_n[8] a_29374_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4973 a_14410_4500# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4974 vcm a_2275_18218# a_5978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4975 vcm a_2275_18218# a_16018_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4976 a_11910_2130# a_2275_2154# a_12002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4977 VSS row_n[14] a_28370_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4978 a_32386_14218# rowon_n[12] a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4979 a_20034_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4980 VDD rowon_n[10] a_27974_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4981 a_8990_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4982 VSS row_n[3] a_23350_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4983 a_10998_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4984 a_33086_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4985 a_27974_1126# a_2275_1150# a_28066_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4986 a_20946_14178# a_2275_14202# a_21038_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4987 a_33998_13174# a_2275_13198# a_34090_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4988 a_4882_8154# a_2275_8178# a_4974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4989 a_5886_4138# a_2275_4162# a_5978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4990 VDD VDD a_26970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4991 a_4974_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4992 a_15014_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4993 a_25454_8516# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4994 VDD rowon_n[6] a_35002_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4995 a_2161_17214# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4996 a_23446_3496# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4997 a_22954_14178# row_n[12] a_23446_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4998 a_8290_10202# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4999 a_18330_10202# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5000 vcm a_2275_10186# a_23046_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5001 a_32386_9198# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5002 VSS row_n[5] a_27366_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5003 VSS row_n[1] a_28370_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5004 a_6982_12170# a_2475_12194# a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5005 a_9902_12170# a_2275_12194# a_9994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5006 a_17022_12170# a_2475_12194# a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5007 VSS row_n[4] a_6282_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5008 a_1957_3158# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5009 a_17326_16226# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5010 vcm a_2275_16210# a_22042_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5011 VSS row_n[7] a_18330_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5012 a_16018_18194# a_2475_18218# a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5013 a_7286_16226# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5014 a_2161_1150# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5015 a_2966_4138# a_2475_4162# a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5016 a_5978_18194# a_2475_18218# a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5017 a_7382_12532# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5018 a_17422_12532# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5019 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5020 a_13310_3174# rowon_n[1] a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5021 vcm a_2275_7174# a_20034_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5022 a_28466_1488# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5023 a_31078_3134# a_2475_3158# a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5024 vcm a_2275_3158# a_21038_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5025 a_16418_18556# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5026 a_26970_8154# a_2275_8178# a_27062_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5027 a_30074_7150# a_2475_7174# a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5028 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5029 a_6378_18556# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5030 vcm a_2275_9182# a_10998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5031 a_31990_9158# row_n[7] a_32482_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5032 a_22042_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5033 a_18426_9520# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5034 VDD VSS a_12914_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5035 VDD rowon_n[3] a_19942_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5036 a_14922_17190# row_n[15] a_15414_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5037 a_26362_15222# rowon_n[13] a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5038 vcm a_2275_13198# a_15014_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5039 VSS row_n[10] a_23350_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5040 VSS VDD a_32386_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5041 a_4882_17190# row_n[15] a_5374_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5042 vcm a_2275_13198# a_4974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5043 a_6982_6146# a_2475_6170# a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5044 vcm a_2275_1150# a_26058_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5045 VSS row_n[9] a_27366_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5046 vcm a_2275_5166# a_25054_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5047 vcm a_2275_8178# a_2966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5048 vcm a_2275_4162# a_3970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5049 a_35094_5142# a_2475_5166# a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5050 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5051 VDD rowon_n[12] a_21950_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5052 a_32082_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5053 a_17326_10202# rowon_n[8] a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5054 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5055 a_7286_10202# rowon_n[8] a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5056 a_18026_2130# a_2475_2154# a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5057 a_31078_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5058 VDD rowon_n[11] a_25966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5059 a_23446_10524# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5060 a_30986_6146# a_2275_6170# a_31078_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5061 VDD rowon_n[5] a_23958_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5062 a_21342_17230# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5063 a_31990_14178# a_2275_14202# a_32082_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5064 a_25358_16226# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5065 a_28370_9198# rowon_n[7] a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5066 VDD rowon_n[0] a_21950_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5067 a_29982_17190# a_2275_17214# a_30074_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5068 vcm a_2275_6170# a_7986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5069 a_9902_2130# row_n[0] a_10394_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5070 a_8290_18234# VDD a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5071 VSS row_n[13] a_5278_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5072 VSS row_n[13] a_15318_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5073 a_20034_15182# a_2475_15206# a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5074 a_12306_12210# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5075 a_21342_8194# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5076 a_27366_2170# rowon_n[0] a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5077 a_22346_4178# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5078 a_24450_18556# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5079 a_24050_14178# a_2475_14202# a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5080 a_16322_11206# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5081 vcm a_2275_11190# a_21038_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5082 VSS row_n[6] a_31382_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5083 a_5278_5182# rowon_n[3] a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5084 a_15318_2170# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5085 a_20946_15182# row_n[13] a_21438_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5086 VSS row_n[12] a_9294_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5087 a_33998_14178# row_n[12] a_34490_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5088 a_15014_13174# a_2475_13198# a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5089 a_6282_11206# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5090 vcm a_2275_10186# a_34090_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5091 a_17326_8194# rowon_n[6] a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5092 a_35002_8154# a_2275_8178# a_35094_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5093 a_19430_5504# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5094 a_4974_13174# a_2475_13198# a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5095 VDD rowon_n[7] a_27974_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5096 vcm a_2275_2154# a_19030_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5097 VDD rowon_n[3] a_28978_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5098 VDD rowon_n[15] a_3878_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5099 VDD rowon_n[15] a_13918_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5100 a_11398_14540# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5101 VDD rowon_n[6] a_6890_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5102 a_15414_13536# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5103 a_11910_10162# row_n[8] a_12402_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5104 a_20034_2130# a_2475_2154# a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5105 VDD rowon_n[14] a_7894_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5106 a_5374_13536# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5107 a_26058_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5108 a_21950_4138# row_n[2] a_22442_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5109 VDD rowon_n[1] a_4882_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5110 a_26362_6186# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5111 vcm a_2275_18218# a_35094_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5112 a_4274_9198# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5113 a_9294_7190# rowon_n[5] a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5114 a_20338_17230# rowon_n[15] a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5115 a_17022_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5116 a_2874_18194# VDD a_3366_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5117 a_12914_18194# VDD a_13406_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5118 a_24354_16226# rowon_n[14] a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5119 vcm a_2275_14202# a_2966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5120 vcm a_2275_14202# a_13006_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5121 VSS row_n[11] a_21342_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5122 a_6982_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5123 a_29070_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5124 a_25966_15182# a_2275_15206# a_26058_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5125 a_30074_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5126 a_3878_9158# row_n[7] a_4370_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5127 a_14010_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5128 a_20946_1126# a_2275_1150# a_21038_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5129 a_19942_5142# a_2275_5166# a_20034_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5130 VDD rowon_n[13] a_19942_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5131 a_5278_11206# rowon_n[9] a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5132 a_15318_11206# rowon_n[9] a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5133 a_16930_8154# row_n[6] a_17422_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5134 a_31078_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5135 a_30074_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5136 a_9994_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5137 a_20338_12210# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5138 a_21438_11528# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5139 a_30378_4178# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5140 a_18330_4178# rowon_n[2] a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5141 a_13006_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5142 a_32386_17230# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5143 a_29070_2130# a_2475_2154# a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5144 VSS row_n[8] a_14314_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5145 vcm a_2275_8178# a_33086_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5146 a_19334_7190# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5147 vcm a_2275_4162# a_34090_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5148 a_4882_11166# a_2275_11190# a_4974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5149 a_14922_11166# a_2275_11190# a_15014_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5150 VSS row_n[8] a_4274_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5151 VSS row_n[5] a_20338_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5152 VSS row_n[1] a_21342_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5153 a_6982_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5154 VSS row_n[14] a_13310_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5155 a_19942_10162# row_n[8] a_20434_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5156 a_8898_7150# row_n[5] a_9390_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5157 a_30378_7190# rowon_n[5] a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5158 a_24962_3134# a_2275_3158# a_25054_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5159 vcm a_2275_17214# a_27062_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5160 VSS row_n[14] a_3270_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5161 a_31078_15182# a_2475_15206# a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5162 VSS row_n[7] a_11302_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5163 a_34090_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5164 a_2874_6146# a_2275_6170# a_2966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5165 a_35094_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5166 VDD rowon_n[10] a_12914_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5167 a_23446_6508# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5168 a_6890_2130# row_n[0] a_7382_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5169 a_29982_4138# row_n[2] a_30474_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5170 VDD rowon_n[2] a_17934_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5171 a_35494_18556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5172 a_31990_15182# row_n[13] a_32482_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5173 a_13006_14178# a_2475_14202# a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5174 a_35094_14178# a_2475_14202# a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5175 VDD rowon_n[10] a_2874_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5176 vcm a_2275_11190# a_32082_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5177 a_14922_9158# a_2275_9182# a_15014_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5178 a_7894_18194# a_2275_18218# a_7986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5179 VDD VDD a_11910_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5180 a_17934_18194# a_2275_18218# a_18026_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5181 a_2966_14178# a_2475_14202# a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5182 a_2161_11190# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5183 VDD a_2161_2154# a_2275_2154# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.615 as=0.342 ps=2.97 w=1.2 l=0.15
X5184 a_21438_1488# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5185 a_13918_2130# a_2275_2154# a_14010_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5186 VSS VDD a_26362_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5187 VSS row_n[3] a_25358_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5188 a_11398_9520# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5189 VSS row_n[6] a_3270_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5190 a_35398_5182# rowon_n[3] a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5191 a_18330_17230# rowon_n[15] a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5192 a_7894_4138# a_2275_4162# a_7986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5193 a_27462_8516# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5194 VSS row_n[11] a_19334_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5195 a_23350_11206# rowon_n[9] a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5196 a_12002_9158# a_2475_9182# a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5197 a_11302_1166# VSS a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5198 a_4974_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5199 a_15014_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5200 a_25454_3496# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5201 a_35398_16226# rowon_n[14] a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5202 VDD rowon_n[1] a_35002_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5203 VDD rowon_n[13] a_17934_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5204 a_10998_2130# a_2475_2154# a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5205 a_8990_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5206 a_34394_9198# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5207 a_16418_7512# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5208 VSS row_n[5] a_29374_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5209 VSS row_n[4] a_8290_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5210 a_23958_16186# a_2275_16210# a_24050_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5211 a_19430_11528# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5212 a_7986_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5213 a_18026_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5214 VSS row_n[13] a_34394_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5215 a_31382_12210# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5216 a_21342_9198# rowon_n[7] a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5217 a_3970_8154# a_2475_8178# a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5218 a_2161_5166# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5219 a_4974_4138# a_2475_4162# a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5220 vcm a_2275_3158# a_23046_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5221 a_11302_15222# rowon_n[13] a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5222 a_35398_11206# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5223 a_28978_8154# a_2275_8178# a_29070_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5224 a_32082_7150# a_2475_7174# a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5225 a_33086_3134# a_2475_3158# a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5226 vcm a_2275_9182# a_13006_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5227 a_20338_2170# rowon_n[0] a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5228 VDD rowon_n[15] a_32994_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5229 a_29070_15182# a_2475_15206# a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5230 a_30474_14540# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5231 vcm a_2275_12194# a_26058_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5232 VSS row_n[9] a_12306_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5233 a_30074_10162# a_2475_10186# a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5234 a_33998_9158# row_n[7] a_34490_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5235 a_24050_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5236 a_34490_13536# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5237 a_30986_10162# row_n[8] a_31478_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5238 a_10298_8194# rowon_n[6] a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5239 VDD rowon_n[3] a_21950_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5240 VDD rowon_n[7] a_20946_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5241 a_9902_5142# row_n[3] a_10394_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5242 vcm a_2275_2154# a_12002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5243 VDD rowon_n[11] a_10906_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5244 a_8990_6146# a_2475_6170# a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5245 vcm a_2275_1150# a_28066_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5246 vcm a_2275_8178# a_4974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5247 vcm a_2275_4162# a_5978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5248 a_10298_16226# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5249 a_2475_3158# a_1957_3158# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X5250 a_32994_6146# a_2275_6170# a_33086_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5251 a_15318_6186# rowon_n[4] a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5252 a_29374_17230# rowon_n[15] a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5253 vcm a_2275_15206# a_18026_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5254 VDD rowon_n[5] a_25966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5255 vcm a_2275_15206# a_7986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5256 a_30378_12210# rowon_n[10] a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5257 VDD rowon_n[4] a_4882_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5258 a_34394_11206# rowon_n[9] a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5259 a_27366_10202# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5260 VDD rowon_n[0] a_23958_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5261 a_22042_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5262 VSS row_n[0] a_19334_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5263 a_24354_4178# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5264 a_23350_8194# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5265 VSS row_n[6] a_33390_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5266 a_29374_2170# rowon_n[0] a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5267 VDD rowon_n[13] a_28978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5268 a_17022_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5269 a_26458_12532# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5270 VDD rowon_n[8] a_29982_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5271 a_7286_5182# rowon_n[3] a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5272 a_6982_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5273 vcm a_2275_8178# a_27062_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5274 VDD rowon_n[6] a_8898_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5275 a_22042_2130# a_2475_2154# a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5276 a_28370_18234# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5277 VSS row_n[14] a_32386_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5278 a_12306_7190# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5279 a_28066_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5280 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5281 VDD rowon_n[1] a_6890_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5282 a_23958_4138# row_n[2] a_24450_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5283 VSS row_n[15] a_8290_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5284 VSS row_n[15] a_18330_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5285 a_23046_17190# a_2475_17214# a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5286 a_27062_16186# a_2475_16210# a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5287 vcm a_2275_13198# a_24050_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5288 a_28370_6186# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5289 VDD VDD a_30986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5290 a_23958_17190# row_n[15] a_24450_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5291 a_18026_15182# a_2475_15206# a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5292 a_9294_13214# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5293 a_19334_13214# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5294 a_6282_9198# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5295 a_27974_16186# row_n[14] a_28466_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5296 a_7986_15182# a_2475_15206# a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5297 a_10906_15182# a_2275_15206# a_10998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5298 a_14922_14178# a_2275_14202# a_15014_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5299 a_4882_14178# a_2275_14202# a_4974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5300 a_8386_15544# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5301 a_18426_15544# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5302 vcm a_2275_6170# a_31078_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5303 a_17326_5182# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5304 a_18938_11166# row_n[9] a_19430_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5305 a_8898_11166# row_n[9] a_9390_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5306 a_5886_9158# row_n[7] a_6378_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5307 a_3970_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5308 a_6890_5142# row_n[3] a_7382_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5309 a_18938_8154# row_n[6] a_19430_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5310 a_22954_1126# a_2275_1150# a_23046_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5311 a_33086_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5312 a_2161_14202# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5313 a_32082_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5314 vcm a_2275_17214# a_12002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5315 a_28370_12210# rowon_n[10] a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5316 a_25966_10162# a_2275_10186# a_26058_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5317 a_20434_8516# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5318 VDD rowon_n[6] a_29982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5319 a_15014_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5320 a_16930_3134# row_n[1] a_17422_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5321 a_27366_18234# VDD a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5322 vcm a_2275_16210# a_5978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5323 vcm a_2275_16210# a_16018_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5324 vcm a_2275_8178# a_35094_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5325 VSS row_n[12] a_28370_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5326 a_28978_17190# a_2275_17214# a_29070_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5327 a_20034_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5328 VDD rowon_n[8] a_27974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5329 VSS row_n[5] a_22346_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5330 VSS row_n[1] a_23350_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5331 a_8990_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5332 a_10998_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5333 a_33086_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5334 a_32386_7190# rowon_n[5] a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5335 VSS row_n[7] a_13310_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5336 a_19030_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5337 a_26058_7150# a_2475_7174# a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5338 a_4882_6146# a_2275_6170# a_4974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5339 VDD rowon_n[14] a_26970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5340 a_4974_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5341 a_15014_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5342 a_25454_6508# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5343 a_8898_2130# row_n[0] a_9390_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5344 VDD rowon_n[4] a_35002_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5345 a_2161_15206# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5346 a_23446_1488# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5347 VSS row_n[10] a_17326_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5348 a_22042_12170# a_2475_12194# a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5349 a_21950_8154# a_2275_8178# a_22042_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5350 a_15926_2130# a_2275_2154# a_16018_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5351 VSS row_n[10] a_7286_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5352 VSS VDD a_16322_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5353 a_21038_18194# a_2475_18218# a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5354 a_22954_12170# row_n[10] a_23446_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5355 VSS VDD a_28370_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5356 VSS row_n[3] a_27366_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5357 VSS VDD a_6282_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5358 a_6982_10162# a_2475_10186# a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5359 a_17022_10162# a_2475_10186# a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5360 a_13406_9520# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5361 VSS row_n[6] a_5278_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5362 a_1957_1150# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5363 VSS row_n[2] a_6282_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5364 a_21950_18194# VDD a_22442_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5365 VDD rowon_n[12] a_15926_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5366 a_17326_14218# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5367 vcm a_2275_14202# a_22042_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5368 a_1957_17214# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5369 a_16018_16186# a_2475_16210# a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5370 VDD rowon_n[12] a_5886_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5371 a_7286_14218# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5372 a_29470_8516# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5373 a_5978_16186# a_2475_16210# a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5374 a_7382_10524# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5375 a_17422_10524# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5376 a_13310_1166# VSS a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5377 vcm a_2275_1150# a_21038_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5378 a_15318_17230# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5379 vcm a_2275_17214# a_20034_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5380 a_14010_9158# a_2475_9182# a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5381 a_31078_1126# a_2475_1150# a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5382 vcm a_2275_5166# a_20034_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5383 a_5278_17230# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5384 a_16418_16548# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5385 a_26970_6146# a_2275_6170# a_27062_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5386 a_27462_3496# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5387 a_30074_5142# a_2475_5166# a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5388 a_6378_16548# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5389 a_31990_7150# row_n[5] a_32482_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5390 a_6378_4500# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5391 a_13006_2130# a_2475_2154# a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5392 vcm a_2275_12194# a_10998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5393 a_18426_7512# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5394 a_14922_15182# row_n[13] a_15414_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5395 a_26362_13214# rowon_n[11] a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5396 vcm a_2275_11190# a_15014_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5397 VSS row_n[8] a_23350_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5398 a_16418_2492# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5399 a_4882_15182# row_n[13] a_5374_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5400 vcm a_2275_11190# a_4974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5401 a_23958_11166# a_2275_11190# a_24050_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5402 a_23350_9198# rowon_n[7] a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5403 a_6982_4138# a_2475_4162# a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5404 a_35094_3134# a_2475_3158# a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5405 vcm a_2275_3158# a_25054_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5406 a_1957_18218# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5407 a_34090_7150# a_2475_7174# a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5408 vcm a_2275_6170# a_2966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5409 VDD rowon_n[10] a_21950_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5410 a_27974_12170# a_2275_12194# a_28066_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5411 vcm a_2275_9182# a_15014_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5412 a_22346_2170# rowon_n[0] a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5413 a_10298_2170# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5414 a_26970_18194# a_2275_18218# a_27062_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5415 a_31078_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5416 VDD rowon_n[9] a_25966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5417 a_12306_8194# rowon_n[6] a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5418 a_29982_8154# a_2275_8178# a_30074_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5419 a_30986_4138# a_2275_4162# a_31078_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5420 VDD rowon_n[7] a_22954_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5421 vcm a_2275_2154# a_14010_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5422 VDD rowon_n[3] a_23958_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5423 VSS VDD a_24354_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5424 a_21342_15222# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5425 a_25358_14218# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5426 a_14314_17230# rowon_n[15] a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5427 a_21038_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5428 a_19030_18194# a_2475_18218# a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5429 a_4274_17230# rowon_n[15] a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5430 a_29982_15182# a_2275_15206# a_30074_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5431 vcm a_2275_4162# a_7986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5432 a_20434_17552# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5433 a_8290_16226# rowon_n[14] a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5434 VSS row_n[11] a_5278_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5435 VSS row_n[11] a_15318_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5436 a_20034_13174# a_2475_13198# a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5437 a_33086_12170# a_2475_12194# a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5438 a_12306_10202# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5439 a_21342_6186# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5440 a_24450_16548# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5441 a_20946_13174# row_n[11] a_21438_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5442 a_10998_12170# a_2475_12194# a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5443 a_4274_7190# rowon_n[5] a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5444 VSS row_n[4] a_31382_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5445 a_5278_3174# rowon_n[1] a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5446 a_33998_12170# row_n[10] a_34490_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5447 a_15014_11166# a_2475_11190# a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5448 a_17326_6186# rowon_n[4] a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5449 a_35002_6146# a_2275_6170# a_35094_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5450 a_4974_11166# a_2475_11190# a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5451 VDD rowon_n[5] a_27974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5452 VDD rowon_n[13] a_3878_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5453 VDD rowon_n[13] a_13918_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5454 a_11398_12532# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5455 VDD rowon_n[4] a_6890_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5456 a_15414_11528# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5457 a_5374_11528# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5458 VDD rowon_n[0] a_25966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5459 a_26058_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5460 a_13310_18234# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5461 VDD VSS a_4882_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5462 a_3270_18234# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5463 vcm a_2275_17214# a_31078_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5464 a_25358_8194# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5465 a_26362_4178# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5466 vcm a_2275_16210# a_35094_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5467 a_11910_8154# row_n[6] a_12402_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5468 VSS row_n[6] a_35398_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5469 a_9294_5182# rowon_n[3] a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5470 a_22042_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5471 a_20338_15222# rowon_n[13] a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5472 vcm a_2275_8178# a_29070_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5473 a_2874_16186# row_n[14] a_3366_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5474 a_12914_16186# row_n[14] a_13406_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5475 a_24354_14218# rowon_n[12] a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5476 VSS row_n[9] a_21342_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5477 a_24050_2130# a_2475_2154# a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5478 a_25054_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5479 a_14314_7190# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5480 VDD rowon_n[1] a_8898_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5481 a_25966_4138# row_n[2] a_26458_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5482 a_29070_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5483 a_25966_13174# a_2275_13198# a_26058_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5484 a_3878_7150# row_n[5] a_4370_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5485 a_19942_3134# a_2275_3158# a_20034_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5486 VDD VDD a_18938_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5487 VDD rowon_n[11] a_19942_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5488 a_8290_9198# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5489 a_16930_6146# row_n[4] a_17422_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5490 a_30074_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5491 a_9994_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5492 a_20338_10202# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5493 a_2475_12194# a_1957_12194# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X5494 a_9902_9158# a_2275_9182# a_9994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5495 a_13310_12210# rowon_n[10] a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5496 a_32386_15222# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5497 a_3270_12210# rowon_n[10] a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5498 a_10906_10162# a_2275_10186# a_10998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5499 a_7286_2170# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5500 vcm a_2275_6170# a_33086_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5501 a_19334_5182# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5502 a_12306_18234# VDD a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5503 VSS VDD a_21342_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5504 VSS row_n[3] a_20338_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5505 VSS row_n[12] a_13310_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5506 a_7894_9158# row_n[7] a_8386_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5507 a_8898_5142# row_n[3] a_9390_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5508 a_24962_1126# a_2275_1150# a_25054_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5509 a_30378_5182# rowon_n[3] a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5510 a_31478_17552# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5511 vcm a_2275_15206# a_27062_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5512 VSS row_n[12] a_3270_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5513 a_31078_13174# a_2475_13198# a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5514 a_35094_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5515 a_2874_4138# a_2275_4162# a_2966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5516 a_34090_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5517 a_3878_17190# a_2275_17214# a_3970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5518 a_13918_17190# a_2275_17214# a_14010_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5519 VDD rowon_n[8] a_12914_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5520 a_22442_8516# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5521 a_35494_16548# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5522 a_31990_13174# row_n[11] a_32482_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5523 VDD rowon_n[8] a_2874_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5524 VDD rowon_n[6] a_31990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5525 a_18938_3134# row_n[1] a_19430_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5526 a_7894_16186# a_2275_16210# a_7986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5527 VDD rowon_n[14] a_11910_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5528 a_17934_16186# a_2275_16210# a_18026_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5529 a_17022_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5530 a_20434_3496# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5531 vcm a_2275_12194# a_30074_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5532 VDD rowon_n[1] a_29982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5533 VSS row_n[1] a_25358_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5534 a_11398_7512# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5535 VSS row_n[5] a_24354_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5536 a_34394_7190# rowon_n[5] a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5537 VSS row_n[4] a_3270_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5538 a_35398_3174# rowon_n[1] a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5539 a_18330_15222# rowon_n[13] a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5540 a_20034_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5541 VSS row_n[7] a_15318_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5542 a_28066_7150# a_2475_7174# a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5543 a_27462_6508# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5544 VSS row_n[9] a_19334_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5545 a_10998_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5546 a_33086_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5547 vcm a_2275_18218# a_19030_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5548 a_5978_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5549 vcm a_2275_18218# a_8990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5550 a_24050_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5551 a_23958_8154# a_2275_8178# a_24050_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5552 a_25454_1488# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5553 a_35398_14218# rowon_n[12] a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5554 VDD VSS a_35002_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5555 a_17934_2130# a_2275_2154# a_18026_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5556 a_23046_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5557 VDD rowon_n[11] a_17934_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5558 VSS row_n[3] a_29374_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5559 a_15414_9520# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5560 a_16418_5504# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5561 VSS row_n[2] a_8290_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5562 a_33390_17230# rowon_n[15] a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5563 a_23958_14178# a_2275_14202# a_24050_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5564 VSS row_n[6] a_7286_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5565 a_7986_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5566 a_18026_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5567 VSS row_n[11] a_34394_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5568 a_31382_10202# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5569 a_3970_6146# a_2475_6170# a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5570 a_2161_3158# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5571 vcm a_2275_1150# a_23046_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5572 a_11302_13214# rowon_n[11] a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5573 a_1957_12194# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5574 a_28978_6146# a_2275_6170# a_29070_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5575 a_33086_1126# a_2475_1150# a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5576 a_29470_3496# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5577 a_32082_5142# a_2475_5166# a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5578 a_6890_9158# a_2275_9182# a_6982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5579 a_29470_17552# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5580 VDD rowon_n[13] a_32994_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5581 a_25966_14178# row_n[12] a_26458_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5582 a_29070_13174# a_2475_13198# a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5583 a_30474_12532# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5584 vcm a_2275_10186# a_26058_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5585 a_33998_7150# row_n[5] a_34490_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5586 a_8386_4500# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5587 a_9994_12170# a_2475_12194# a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5588 a_12914_12170# a_2275_12194# a_13006_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5589 a_15014_2130# a_2475_2154# a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5590 a_2874_12170# a_2275_12194# a_2966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5591 a_34490_11528# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5592 a_10298_6186# rowon_n[4] a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5593 a_31990_2130# row_n[0] a_32482_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5594 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5595 a_11910_18194# a_2275_18218# a_12002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5596 VDD rowon_n[9] a_10906_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5597 VDD rowon_n[5] a_20946_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5598 a_18426_2492# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5599 a_8990_4138# a_2475_4162# a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5600 a_19030_9158# a_2475_9182# a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5601 vcm a_2275_6170# a_4974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5602 a_10298_14218# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5603 a_2475_1150# a_1957_1150# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X5604 a_24354_2170# rowon_n[0] a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5605 a_32994_4138# a_2275_4162# a_33086_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5606 a_14314_8194# rowon_n[6] a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5607 vcm a_2275_8178# a_22042_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5608 a_15318_4178# rowon_n[2] a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5609 a_17934_17190# row_n[15] a_18426_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5610 a_29374_15222# rowon_n[13] a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5611 vcm a_2275_13198# a_18026_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5612 VSS row_n[10] a_26362_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5613 vcm a_2275_2154# a_16018_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5614 VDD rowon_n[3] a_25966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5615 a_7894_17190# row_n[15] a_8386_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5616 vcm a_2275_13198# a_7986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5617 a_31078_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5618 a_30378_10202# rowon_n[8] a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5619 VDD rowon_n[6] a_3878_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5620 a_22042_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5621 a_23046_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5622 VDD rowon_n[12] a_24962_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5623 a_13006_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5624 a_35094_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5625 a_2966_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5626 a_23350_6186# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5627 VSS row_n[4] a_33390_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5628 VDD rowon_n[2] a_14922_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5629 VDD rowon_n[11] a_28978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5630 a_26458_10524# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5631 a_29982_10162# a_2275_10186# a_30074_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5632 a_6282_7190# rowon_n[5] a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5633 a_7286_3174# rowon_n[1] a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5634 vcm a_2275_6170# a_27062_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5635 a_31382_18234# VDD a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5636 a_24354_17230# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5637 VDD rowon_n[4] a_8898_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5638 a_28370_16226# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5639 VSS row_n[12] a_32386_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5640 a_12306_5182# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5641 VDD rowon_n[0] a_27974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5642 a_28066_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5643 a_19942_18194# a_2275_18218# a_20034_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5644 a_32994_17190# a_2275_17214# a_33086_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5645 VDD VSS a_6890_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5646 VSS row_n[13] a_8290_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5647 VSS row_n[13] a_18330_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5648 a_23046_15182# a_2475_15206# a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5649 a_27062_14178# a_2475_14202# a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5650 a_19334_11206# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5651 vcm a_2275_11190# a_24050_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5652 a_13918_8154# row_n[6] a_14410_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5653 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5654 a_28370_4178# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5655 a_27462_18556# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5656 VDD rowon_n[14] a_30986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5657 a_23958_15182# row_n[13] a_24450_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5658 a_18026_13174# a_2475_13198# a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5659 a_9294_11206# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5660 a_7986_13174# a_2475_13198# a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5661 a_10906_13174# a_2275_13198# a_10998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5662 VDD rowon_n[15] a_6890_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5663 VDD rowon_n[15] a_16930_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5664 a_11910_3134# row_n[1] a_12402_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5665 a_18426_13536# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5666 a_8386_13536# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5667 vcm a_2275_8178# a_30074_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5668 a_16322_7190# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5669 a_17326_3174# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5670 vcm a_2275_4162# a_31078_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5671 a_27974_4138# row_n[2] a_28466_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5672 a_5886_7150# row_n[5] a_6378_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5673 a_3970_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5674 a_18938_6146# row_n[4] a_19430_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5675 a_21038_7150# a_2475_7174# a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5676 a_32082_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5677 vcm a_2275_15206# a_12002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5678 a_29070_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5679 a_28370_10202# rowon_n[8] a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5680 a_20434_6508# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5681 a_3878_2130# row_n[0] a_4370_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5682 VDD rowon_n[4] a_29982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5683 a_16930_1126# VDD a_17422_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5684 a_15926_18194# VDD a_16418_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5685 a_27366_16226# rowon_n[14] a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5686 vcm a_2275_14202# a_5978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5687 vcm a_2275_14202# a_16018_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5688 a_9994_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5689 a_9294_2170# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5690 a_5886_18194# VDD a_6378_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5691 vcm a_2275_6170# a_35094_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5692 a_10906_2130# a_2275_2154# a_10998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5693 a_28978_15182# a_2275_15206# a_29070_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5694 a_20034_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5695 VSS VDD a_23350_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5696 VSS row_n[3] a_22346_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5697 a_10998_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5698 a_33086_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5699 a_32386_5182# rowon_n[3] a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5700 a_23350_12210# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5701 a_4882_4138# a_2275_4162# a_4974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5702 a_26058_5142# a_2475_5166# a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5703 a_24450_8516# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5704 a_22346_18234# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5705 VDD rowon_n[6] a_33998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5706 a_2161_13198# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5707 a_22442_14540# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5708 VSS row_n[8] a_17326_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5709 a_22042_10162# a_2475_10186# a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5710 VSS a_2161_8178# a_2275_8178# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X5711 a_21950_6146# a_2275_6170# a_22042_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5712 VDD rowon_n[1] a_31990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5713 a_22442_3496# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5714 a_7894_11166# a_2275_11190# a_7986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5715 a_17934_11166# a_2275_11190# a_18026_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5716 VSS row_n[8] a_7286_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5717 a_30986_18194# a_2275_18218# a_31078_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5718 VSS row_n[14] a_16322_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5719 a_21038_16186# a_2475_16210# a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5720 a_22954_10162# row_n[8] a_23446_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5721 VSS row_n[1] a_27366_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5722 VSS row_n[14] a_6282_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5723 a_19334_9198# rowon_n[7] a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5724 a_31382_9198# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5725 a_13406_7512# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5726 VSS row_n[4] a_5278_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5727 a_21950_16186# row_n[14] a_22442_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5728 VDD rowon_n[10] a_15926_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5729 VSS row_n[7] a_17326_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5730 a_1957_15206# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5731 a_16018_14178# a_2475_14202# a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5732 VDD rowon_n[10] a_5886_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5733 a_29470_6508# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5734 a_11398_2492# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5735 VDD VDD a_14922_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5736 a_5978_14178# a_2475_14202# a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5737 VDD VDD a_4882_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5738 a_15318_15222# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5739 vcm a_2275_15206# a_20034_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5740 a_7986_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5741 VSS row_n[0] a_16322_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5742 a_30074_3134# a_2475_3158# a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5743 vcm a_2275_3158# a_20034_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5744 a_14010_17190# a_2475_17214# a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5745 a_5278_15222# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5746 a_25966_8154# a_2275_8178# a_26058_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5747 a_27462_1488# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5748 a_26970_4138# a_2275_4162# a_27062_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5749 a_3970_17190# a_2475_17214# a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5750 vcm a_2275_9182# a_9994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5751 VDD rowon_n[7] a_18938_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5752 a_30986_9158# row_n[7] a_31478_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5753 a_31990_5142# row_n[3] a_32482_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5754 a_14410_17552# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5755 a_10906_14178# row_n[12] a_11398_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5756 vcm a_2275_10186# a_10998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5757 a_17422_9520# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5758 VSS row_n[6] a_9294_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5759 a_18426_5504# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5760 a_4370_17552# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5761 a_22346_12210# rowon_n[10] a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5762 a_14922_13174# row_n[11] a_15414_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5763 a_26362_11206# rowon_n[9] a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5764 a_4882_13174# row_n[11] a_5374_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5765 a_18026_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5766 vcm a_2275_1150# a_25054_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5767 a_35094_1126# a_2475_1150# a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5768 a_1957_16210# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5769 a_7986_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5770 a_1957_6170# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5771 vcm a_2275_4162# a_2966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5772 a_34090_5142# a_2475_5166# a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5773 VDD rowon_n[8] a_21950_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5774 a_8898_9158# a_2275_9182# a_8990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5775 a_17022_2130# a_2475_2154# a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5776 VSS row_n[15] a_20338_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5777 a_26970_16186# a_2275_16210# a_27062_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5778 a_31078_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5779 a_12306_6186# rowon_n[4] a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5780 a_29982_6146# a_2275_6170# a_30074_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5781 VDD rowon_n[5] a_22954_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5782 a_33998_2130# row_n[0] a_34490_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5783 VSS row_n[14] a_24354_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5784 a_21342_13214# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5785 a_34394_12210# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5786 a_14314_15222# rowon_n[13] a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5787 VSS row_n[10] a_11302_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5788 VDD rowon_n[0] a_20946_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5789 a_21038_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5790 a_19030_16186# a_2475_16210# a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5791 a_4274_15222# rowon_n[13] a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5792 a_29982_13174# a_2275_13198# a_30074_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5793 VDD VDD a_22954_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5794 a_20434_15544# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5795 a_8290_14218# rowon_n[12] a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5796 a_33486_14540# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5797 vcm a_2275_12194# a_29070_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5798 VSS row_n[9] a_5278_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5799 VSS row_n[9] a_15318_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5800 a_20034_11166# a_2475_11190# a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5801 a_33086_10162# a_2475_10186# a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5802 a_20338_8194# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5803 a_26362_2170# rowon_n[0] a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5804 a_21342_4178# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5805 a_20946_11166# row_n[9] a_21438_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5806 a_10998_10162# a_2475_10186# a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5807 a_5978_9158# a_2475_9182# a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5808 VSS row_n[6] a_30378_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5809 a_4274_5182# rowon_n[3] a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5810 a_5278_1166# VSS a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5811 VSS row_n[2] a_31382_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5812 VDD rowon_n[12] a_9902_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5813 a_33998_10162# row_n[8] a_34490_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5814 a_35002_4138# a_2275_4162# a_35094_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5815 a_17326_4178# rowon_n[2] a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5816 a_16322_8194# rowon_n[6] a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5817 vcm a_2275_8178# a_24050_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5818 vcm a_2275_2154# a_18026_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5819 VDD rowon_n[3] a_27974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5820 VDD rowon_n[11] a_3878_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5821 VDD rowon_n[11] a_13918_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5822 a_11398_10524# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5823 VDD rowon_n[6] a_5886_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5824 a_25054_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5825 a_26058_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5826 a_13310_16226# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5827 VDD rowon_n[1] a_3878_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5828 a_31478_4500# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5829 a_20946_4138# row_n[2] a_21438_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5830 a_12002_18194# a_2475_18218# a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5831 a_34090_18194# a_2475_18218# a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5832 a_3270_16226# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5833 vcm a_2275_15206# a_31078_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5834 a_25358_6186# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5835 a_35002_18194# VDD a_35494_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5836 vcm a_2275_14202# a_35094_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5837 a_3270_9198# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5838 a_11910_6146# row_n[4] a_12402_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5839 VSS row_n[4] a_35398_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5840 a_9294_3174# rowon_n[1] a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5841 VDD rowon_n[2] a_16930_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5842 a_8290_7190# rowon_n[5] a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5843 a_12402_18556# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5844 a_19334_18234# VDD a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5845 a_20338_13214# rowon_n[11] a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5846 vcm a_2275_6170# a_29070_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5847 vcm a_2275_9182# a_6982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5848 a_25054_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5849 a_21950_12170# a_2275_12194# a_22042_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5850 a_14314_5182# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5851 VDD VSS a_8898_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5852 a_29070_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5853 a_2874_9158# row_n[7] a_3366_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5854 a_3878_5142# row_n[3] a_4370_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5855 a_19942_1126# a_2275_1150# a_20034_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5856 VDD rowon_n[14] a_18938_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5857 VDD rowon_n[9] a_19942_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5858 a_15926_8154# row_n[6] a_16418_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5859 a_30074_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5860 a_9994_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5861 VSS row_n[15] a_31382_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5862 a_2475_10186# a_1957_10186# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.615 w=1.2 l=0.15
X5863 a_13918_3134# row_n[1] a_14410_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5864 a_13310_10202# rowon_n[8] a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5865 a_12002_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5866 VSS row_n[14] a_35398_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5867 a_32386_13214# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5868 a_3270_10202# rowon_n[8] a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5869 a_18330_7190# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5870 a_19334_3174# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5871 vcm a_2275_4162# a_33086_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5872 a_26058_17190# a_2475_17214# a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5873 a_12306_16226# rowon_n[14] a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5874 VSS row_n[1] a_20338_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5875 a_7894_7150# row_n[5] a_8386_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5876 a_30378_3174# rowon_n[1] a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5877 VDD VDD a_33998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5878 a_26970_17190# row_n[15] a_27462_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5879 a_31478_15544# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5880 vcm a_2275_13198# a_27062_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5881 a_31078_11166# a_2475_11190# a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5882 a_34090_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5883 a_3878_15182# a_2275_15206# a_3970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5884 a_13918_15182# a_2275_15206# a_14010_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5885 VSS row_n[7] a_10298_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5886 a_23046_7150# a_2475_7174# a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5887 a_22442_6508# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5888 a_5886_2130# row_n[0] a_6378_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5889 a_17934_14178# a_2275_14202# a_18026_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5890 a_31990_11166# row_n[9] a_32482_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5891 VDD rowon_n[4] a_31990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5892 a_18938_1126# en_bit_n[2] a_19430_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5893 a_7894_14178# a_2275_14202# a_7986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5894 a_20434_1488# en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5895 a_29982_14178# row_n[12] a_30474_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5896 vcm a_2275_10186# a_30074_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5897 VDD VSS a_29982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5898 a_12914_2130# a_2275_2154# a_13006_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5899 VSS VDD a_25358_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5900 VSS row_n[3] a_24354_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5901 a_10394_9520# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5902 a_11398_5504# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5903 a_35398_1166# VSS a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5904 VSS row_n[2] a_3270_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5905 a_34394_5182# rowon_n[3] a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5906 a_18330_13214# rowon_n[11] a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5907 a_28978_10162# a_2275_10186# a_29070_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5908 a_28066_5142# a_2475_5166# a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5909 vcm a_2275_16210# a_8990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5910 vcm a_2275_16210# a_19030_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5911 a_23958_6146# a_2275_6170# a_24050_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5912 a_24450_3496# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5913 VDD rowon_n[1] a_33998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5914 a_23046_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5915 VDD rowon_n[9] a_17934_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5916 VSS row_n[1] a_29374_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5917 a_3366_4500# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5918 a_33390_9198# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5919 a_15414_7512# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5920 VSS row_n[15] a_29374_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5921 a_33390_15222# rowon_n[13] a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5922 VSS row_n[10] a_30378_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5923 a_16018_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5924 VSS row_n[4] a_7286_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5925 a_7986_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5926 a_18026_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5927 VSS row_n[9] a_34394_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5928 a_32386_2170# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5929 a_2161_1150# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5930 a_13406_2492# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5931 a_3970_4138# a_2475_4162# a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5932 a_9994_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5933 a_25054_12170# a_2475_12194# a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5934 a_11302_11206# rowon_n[9] a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5935 a_1957_10186# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5936 a_27974_8154# a_2275_8178# a_28066_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5937 a_29470_1488# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5938 VSS row_n[0] a_18330_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5939 a_32082_3134# a_2475_3158# a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5940 a_28978_4138# a_2275_4162# a_29070_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5941 a_29470_15544# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5942 VDD rowon_n[11] a_32994_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5943 a_25966_12170# row_n[10] a_26458_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5944 a_29070_11166# a_2475_11190# a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5945 a_30474_10524# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5946 a_32994_9158# row_n[7] a_33486_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5947 a_33998_5142# row_n[3] a_34490_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5948 a_9994_10162# a_2475_10186# a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5949 a_10298_4178# rowon_n[2] a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5950 a_11910_16186# a_2275_16210# a_12002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5951 VDD rowon_n[12] a_8898_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5952 vcm a_2275_2154# a_10998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5953 VDD rowon_n[3] a_20946_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5954 a_16930_7150# a_2275_7174# a_17022_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5955 vcm a_2275_17214# a_23046_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5956 a_8290_17230# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5957 a_18330_17230# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5958 vcm a_2275_4162# a_4974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5959 VDD rowon_n[2] a_9902_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5960 vcm a_2275_12194# a_14010_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5961 vcm a_2275_12194# a_3970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5962 a_14314_6186# rowon_n[4] a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5963 vcm a_2275_6170# a_22042_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5964 a_17934_15182# row_n[13] a_18426_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5965 a_29374_13214# rowon_n[11] a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5966 vcm a_2275_11190# a_18026_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5967 VSS row_n[8] a_26362_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5968 a_7894_15182# row_n[13] a_8386_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5969 vcm a_2275_11190# a_7986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5970 a_26970_11166# a_2275_11190# a_27062_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5971 VDD rowon_n[4] a_3878_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5972 VDD rowon_n[0] a_22954_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5973 a_23046_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5974 VDD rowon_n[10] a_24962_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5975 a_28370_2170# rowon_n[0] a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5976 VSS row_n[2] a_33390_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5977 a_23350_4178# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5978 VDD rowon_n[9] a_28978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5979 a_7986_9158# a_2475_9182# a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5980 VSS row_n[6] a_32386_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5981 a_6282_5182# rowon_n[3] a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5982 a_7286_1166# VSS a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5983 VSS a_2161_18218# a_2275_18218# VSS sky130_fd_pr__nfet_01v8 ad=0.1245 pd=1.015 as=0.171 ps=1.77 w=0.6 l=0.15
X5984 vcm a_2275_8178# a_26058_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5985 vcm a_2275_4162# a_27062_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5986 VSS VDD a_27366_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5987 a_31382_16226# rowon_n[14] a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5988 a_24354_15222# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5989 VDD rowon_n[6] a_7894_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5990 a_2475_6170# a_1957_6170# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.1245 ps=1.015 w=0.6 l=0.15
X5991 a_17326_17230# rowon_n[15] a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5992 a_28370_14218# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5993 a_11302_7190# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5994 a_28066_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5995 a_12306_3174# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5996 a_7286_17230# rowon_n[15] a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5997 a_19942_16186# a_2275_16210# a_20034_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5998 a_32994_15182# a_2275_15206# a_33086_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5999 a_31990_9158# a_2275_9182# a_32082_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6000 a_27062_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6001 a_22954_4138# row_n[2] a_23446_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6002 a_3970_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6003 a_14010_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6004 a_23446_17552# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6005 VSS row_n[11] a_8290_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6006 VSS row_n[11] a_18330_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6007 a_23046_13174# a_2475_13198# a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6008 VDD rowon_n[1] a_5886_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6009 a_33486_4500# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6010 a_13918_6146# row_n[4] a_14410_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6011 a_27462_16548# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6012 a_23958_13174# row_n[11] a_24450_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6013 a_18026_11166# a_2475_11190# a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6014 a_5278_9198# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6015 a_7986_11166# a_2475_11190# a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6016 VDD rowon_n[13] a_6890_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6017 VDD rowon_n[13] a_16930_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6018 vcm a_2275_9182# a_8990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6019 a_11910_1126# VDD a_12402_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6020 a_18426_11528# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6021 a_4274_2170# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6022 a_8386_11528# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6023 vcm a_2275_6170# a_30074_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6024 a_16322_5182# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6025 a_17326_1166# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6026 a_16322_18234# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6027 vcm a_2275_18218# a_21038_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6028 a_6282_18234# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6029 vcm a_2275_17214# a_34090_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6030 a_5886_5142# row_n[3] a_6378_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6031 a_4882_9158# row_n[7] a_5374_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6032 a_17934_8154# row_n[6] a_18426_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6033 a_25054_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6034 a_32082_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6035 a_21038_5142# a_2475_5166# a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6036 a_11910_17190# row_n[15] a_12402_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6037 vcm a_2275_13198# a_12002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6038 a_14010_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6039 a_15926_3134# row_n[1] a_16418_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6040 a_5886_16186# row_n[14] a_6378_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6041 a_15926_16186# row_n[14] a_16418_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6042 a_27366_14218# rowon_n[12] a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6043 a_27366_9198# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6044 vcm a_2275_4162# a_35094_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6045 a_28066_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6046 a_28978_13174# a_2275_13198# a_29070_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6047 VSS row_n[1] a_22346_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6048 a_31382_7190# rowon_n[5] a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6049 a_32386_3174# rowon_n[1] a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6050 a_23350_10202# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6051 VSS row_n[7] a_12306_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6052 a_26058_3134# a_2475_3158# a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6053 a_25054_7150# a_2475_7174# a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6054 a_24450_6508# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6055 a_7894_2130# row_n[0] a_8386_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6056 a_22346_16226# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6057 a_16322_12210# rowon_n[10] a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6058 a_26970_9158# row_n[7] a_27462_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6059 VDD rowon_n[4] a_33998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6060 a_6282_12210# rowon_n[10] a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6061 a_2161_11190# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X6062 a_13918_10162# a_2275_10186# a_14010_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6063 a_2966_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6064 VSS row_n[0] a_11302_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6065 a_22442_12532# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6066 a_3878_10162# a_2275_10186# a_3970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6067 a_20946_8154# a_2275_8178# a_21038_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6068 a_22442_1488# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6069 VDD VSS a_31990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6070 a_21950_4138# a_2275_4162# a_22042_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6071 a_5278_18234# VDD a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6072 a_15318_18234# VDD a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6073 a_31078_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6074 a_14922_2130# a_2275_2154# a_15014_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6075 a_21438_18556# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6076 a_30986_16186# a_2275_16210# a_31078_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6077 VSS row_n[12] a_16322_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6078 a_21038_14178# a_2475_14202# a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6079 VSS VDD a_27366_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6080 VSS row_n[12] a_6282_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6081 a_12402_9520# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6082 VSS row_n[6] a_4274_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6083 a_13406_5504# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6084 VSS row_n[2] a_5278_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6085 a_16930_17190# a_2275_17214# a_17022_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6086 VDD rowon_n[8] a_15926_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6087 a_6890_17190# a_2275_17214# a_6982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6088 VDD rowon_n[8] a_5886_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6089 VSS row_n[15] a_4274_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6090 VSS row_n[15] a_14314_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6091 VDD rowon_n[14] a_14922_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6092 VDD rowon_n[14] a_4882_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6093 a_15318_13214# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6094 vcm a_2275_13198# a_20034_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6095 vcm a_2275_1150# a_20034_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6096 a_30074_1126# a_2475_1150# a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6097 a_19942_17190# row_n[15] a_20434_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6098 a_14010_15182# a_2475_15206# a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6099 a_5278_13214# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6100 vcm a_2275_12194# a_33086_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6101 a_25966_6146# a_2275_6170# a_26058_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 VPWR VGND B1 Y A1 A2 VNB VPB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X3 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15 M=4
X4 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15 M=4
X5 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15 M=4
.ends

.subckt sky130_fd_sc_hd__o211ai_1 VGND VPWR A1 Y C1 B1 A2 VNB VPB
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt adc_inverter in out VDD VSS
X0 out in VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.0651 ps=0.73 w=0.42 l=0.15 M=2
X1 out in VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt adc_nor a b q VDD VSS
X0 a_312_106# b q VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1 VSS b q VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 q a a_120_106# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3 VDD a a_312_106# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4 q a VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5 a_120_106# b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
.ends

.subckt adc_nor_latch qn q s r VDD VSS
X0 a_806_530# qn VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1 q r a_806_530# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2 q r VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3 a_998_530# qn q VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4 VSS qn q VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 VDD r a_998_530# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6 a_480_530# q qn VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X7 qn s VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X8 VSS q qn VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_288_530# q VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X10 qn s a_288_530# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X11 VDD s a_480_530# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
.ends

.subckt adc_noise_decoup_cell2 nmoscap_bot nmoscap_top mimcap_bot mimcap_top pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=5.1 w=18.9
X1 nmoscap_top nmoscap_bot pwell sky130_fd_pr__cap_var_lvt w=18.4 l=3.9
.ends

.subckt adc_comp_buffer out in VDD VSS
X0 out a_26_n216# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15 M=2
X1 VSS a_26_n216# out VSS sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15 M=2
X2 VSS in a_26_n216# VSS sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X3 VDD in a_26_n216# VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
.ends

.subckt adc_comp_circuit bp bn on op a_30_n1001# a_1611_n1292# adc_comp_buffer_0/out
+ a_470_n1001# a_12_n446# VGND adc_comp_buffer_1/out VPWR
Xadc_noise_decoup_cell2_0 VGND op VGND VGND VGND adc_noise_decoup_cell2
Xadc_noise_decoup_cell2_1 VGND on VGND VGND VGND adc_noise_decoup_cell2
Xadc_comp_buffer_0 adc_comp_buffer_0/out bn VPWR VGND adc_comp_buffer
Xadc_comp_buffer_1 adc_comp_buffer_1/out bp VPWR VGND adc_comp_buffer
X0 VPWR a_12_n446# on VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15 M=4
X1 VGND a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15 M=8
X2 bp a_1611_n1292# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.31 ps=2.31 w=2 l=0.15
X3 a_1090_n348# bn VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15 M=2
X4 a_1877_n348# op a_1877_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=2.9 ps=22.9 w=2 l=0.15
X5 op a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15 M=4
X6 VGND bn bp VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7 a_n28_n1170# a_30_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=5.075 pd=43.12 as=0.58 ps=4.58 w=2 l=0.15
X8 op a_30_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15 M=4
X9 on a_470_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15 M=4
X10 a_n28_n1170# a_470_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X11 bp on a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15 M=2
X12 a_1877_n348# bp VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15 M=2
X13 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=55.88 pd=188.82 as=0.62 ps=4.62 w=2 l=0.15 M=2
X14 a_n28_n1170# a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0725 ps=0.79 w=0.5 l=0.15 M=2
X15 bn bp VGND VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X16 a_1877_n348# op bn VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15 M=2
X17 VGND a_1611_n1292# bn VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.31 as=0.33 ps=2.33 w=2 l=0.15
X18 a_1090_n348# bn a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=2.9 pd=22.9 as=0.29 ps=2.29 w=2 l=0.15
X19 a_1090_n348# on a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.15
X20 VPWR a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=2.75003 pd=22.965 as=0.155 ps=1.62 w=0.5 l=0.15 M=2
X21 a_1877_n348# bp a_1877_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt adc_comp_latch clk inp inn comp_trig latch_qn latch_q VDD VSUBS VSS
Xadc_inverter_1 adc_inverter_1/in adc_inverter_1/out VDD VSS adc_inverter
Xadc_inverter_2 clk adc_inverter_1/in VDD VSS adc_inverter
Xadc_nor_0 adc_nor_0/a adc_nor_0/b comp_trig VDD VSS adc_nor
Xadc_nor_latch_0 latch_qn latch_q adc_nor_0/b adc_nor_0/a VDD VSS adc_nor_latch
Xadc_comp_circuit_0 adc_comp_circuit_0/bp adc_comp_circuit_0/bn adc_comp_circuit_0/on
+ adc_comp_circuit_0/op inn adc_inverter_1/in adc_nor_0/a inp adc_inverter_1/out VSS
+ adc_nor_0/b VDD adc_comp_circuit
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR X A1 A2 B1 C1 VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR X D C B A_N VNB VPB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPWR VGND A1 B1_N Y A2 VNB VPB
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 VGND VPWR A1 A2 B2 B1 X VNB VPB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15 M=2
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X6 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X7 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X9 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 VGND VPWR X B1 A2 A1 VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15 M=2
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15 M=2
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND X A B VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15 M=2
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X3 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 VPWR VGND C1 B2 B1 A1 A2 X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15 M=2
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VPWR VGND X A1_N A2_N B2 B1 VNB VPB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X C1 A2 A1 B1 VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt scboundary VDD VSS
X0 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.2484 pd=2.1 as=0.4761 ps=4.14 w=0.69 l=0.71
.ends

.subckt sky130_fd_sc_hd__nand2_4 VGND VPWR B Y A VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=4
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=4
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
.ends

.subckt sky130_fd_sc_hd__o31a_1 VGND VPWR X A1 A2 A3 B1 VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND Q SET_B D CLK VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 VGND VPWR A2 B1 Y A1 VNB VPB
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15 M=4
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15 M=4
X3 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X4 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15 M=4
X5 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15 M=4
.ends

.subckt sky130_mm_sc_hd_dlyPoly5ns VPWR VGND in out mid VNB VPB
X0 a_1691_329# out VGND VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=2.2 as=0.132 ps=1.13 w=0.8 l=0.15 M=2
X1 a_1691_329# mid VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.13 as=0.24 ps=2.2 w=0.8 l=0.15
X2 out mid a_1691_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=2.2 as=0.132 ps=1.13 w=0.8 l=0.15
X3 VGND mid VGND VNB sky130_fd_pr__nfet_01v8 ad=1.0453 pd=9.52 as=0.39875 ps=3.33 w=1.375 l=2.045
X4 a_1632_71# mid VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.126 ps=1.44 w=0.42 l=0.15
X5 VPWR out a_1632_71# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15 M=2
X6 out mid a_1632_71# VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 mid in VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.232 pd=2.18 as=0.232 ps=2.18 w=0.8 l=1.42
X8 mid in VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=3.69
.ends

.subckt sky130_fd_sc_hd__nor2b_1 VGND VPWR B_N A Y VNB VPB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1573 pd=1.39 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.1573 ps=1.39 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__bufbuf_8 VGND VPWR A X VNB VPB
X0 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=3
X1 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=8
X2 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=8
X3 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15 M=3
X4 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5 a_206_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt adc_clkgen_with_edgedetect VDD clk_comp_out clk_dig_out dlycontrol1_in[0]
+ dlycontrol1_in[1] dlycontrol1_in[2] dlycontrol1_in[3] dlycontrol1_in[4] dlycontrol2_in[0]
+ dlycontrol2_in[1] dlycontrol2_in[2] dlycontrol2_in[3] dlycontrol2_in[4] dlycontrol3_in[0]
+ dlycontrol3_in[1] dlycontrol3_in[2] dlycontrol3_in[3] dlycontrol3_in[4] dlycontrol4_in[0]
+ dlycontrol4_in[1] dlycontrol4_in[2] dlycontrol4_in[3] dlycontrol4_in[4] dlycontrol4_in[5]
+ ena_in enable_dlycontrol_in ndecision_finish_in sample_n_in sample_n_out sample_p_in
+ sample_p_out start_conv_in VSS VSUBS
XFILLER_10_317 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[0\]
+ dlycontrol2_in[0] VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_10_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A dlycontrol1_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.clk_dig_delayed_w
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_14_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.or1 VSS VDD clkgen.enable_loop_in edgedetect.start_conv_edge_w edgedetect.ena_in
+ VSS VDD sky130_fd_sc_hd__or2_1
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_334 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[1\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[1\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_3_271 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A dlycontrol2_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[2\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[3\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[4\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_5_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A dlycontrol3_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[1\]
+ dlycontrol4_in[1] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_283 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_198 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_304 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_B edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit_in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.nor1 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out
+ edgedetect.start_conv_edge_w VSS VDD sky130_fd_sc_hd__nor2b_1
XFILLER_7_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.or1_A edgedetect.start_conv_edge_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xdelay_sample_p11 VDD VSS sample_p_in sample_p_1 delay_sample_p11/mid VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_295 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[1\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[1\]
+ dlycontrol3_in[1] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_0_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_265 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_302 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_2_316 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.or1_B edgedetect.ena_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_167 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_328 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.nor1 VSS VDD clkgen.enable_loop_in clkgen.clk_dig_delayed_w clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ VSS VDD sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_B clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[2\]
+ dlycontrol1_in[2] VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_14_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A dlycontrol1_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_inbuf_3_A ndecision_finish_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.clkdig_inverter VDD VSS clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out
+ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_232 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_320 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A dlycontrol2_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_315 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_304 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_277 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xdelay_sample_n12 VDD VSS sample_n_in sample_n_1 delay_sample_n12/mid VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_7_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinbuf_1 VSS VDD edgedetect.ena_in ena_in VSS VDD sky130_fd_sc_hd__buf_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[3\]
+ dlycontrol2_in[3] VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[2\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[2\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_19_327 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[3\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XPHY_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[4\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_8_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinbuf_2 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in start_conv_in VSS
+ VDD sky130_fd_sc_hd__buf_1
XFILLER_12_152 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_9_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_inbuf_1_A ena_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xinbuf_3 VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in ndecision_finish_in
+ VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_16_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_164 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A dlycontrol4_in[5] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[4\]
+ dlycontrol4_in[4] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_1_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B clkgen.clk_dig_out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_284 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[0\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_2_280 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_306 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_1_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[4\]
+ dlycontrol3_in[4] VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_1_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_242 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A dlycontrol1_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_292 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_314 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_290 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[0\]
+ dlycontrol1_in[0] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_12_326 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XPHY_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XPHY_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_244 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_2_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.enablebuffer VDD VSS edgedetect.dly_315ns_1.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_18_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_302 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_195 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A dlycontrol4_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.enablebuffer VDD VSS clkgen.delay_155ns_1.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[3\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[3\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_13_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[1\]
+ dlycontrol2_in[1] VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_312 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_304 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[4\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_2_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_314 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_292 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_324 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_10_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_308 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A1 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_326 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[2\]
+ dlycontrol4_in[2] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_1_307 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[0\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_5_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_336 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[1\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_2_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A dlycontrol3_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.clk_dig_out VSS VDD
+ VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[2\]
+ dlycontrol3_in[2] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_B clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_0_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_285 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_244 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A dlycontrol4_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[3\]
+ dlycontrol1_in[3] VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_10_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_318 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_298 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[4\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_0_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A dlycontrol2_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_278 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.enablebuffer VDD VSS clkgen.delay_155ns_2.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_2_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A dlycontrol3_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[4\]
+ dlycontrol2_in[4] VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_8_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_A1 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_291 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_290 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_271 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_315 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[0\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[0\]
+ dlycontrol4_in[0] VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[0\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[1\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[2\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[5\]
+ dlycontrol4_in[5] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_2_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_283 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_327 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_11_179 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_44 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_A1 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_304 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[0\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[0\]
+ dlycontrol3_in[0] VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_A0 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A dlycontrol4_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_295 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_339 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_inbuf_2_A start_conv_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_3_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutbuf_1 VSS VDD clkgen.clk_dig_out clk_dig_out VSS VDD sky130_fd_sc_hd__bufbuf_8
XFILLER_14_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit_in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A dlycontrol1_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[1\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[1\]
+ dlycontrol1_in[1] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_15_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_edgedetect.nor1_B_N edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A dlycontrol2_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_198 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_2 VSS VDD clkgen.clk_comp_out clk_comp_out VSS VDD sky130_fd_sc_hd__bufbuf_8
XFILLER_6_334 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A dlycontrol3_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_262 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_306 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutbuf_3 VSS VDD sample_p_1 sample_p_out VSS VDD sky130_fd_sc_hd__bufbuf_8
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_14_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_outbuf_1_A clkgen.clk_dig_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_9_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_195 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.clk_comp_out
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[5\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[5\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_6_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutbuf_4 VSS VDD sample_n_1 sample_n_out VSS VDD sky130_fd_sc_hd__bufbuf_8
Xclkgen.delay_155ns_3.enablebuffer VDD VSS clkgen.delay_155ns_3.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[2\]
+ dlycontrol2_in[2] VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_298 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_257 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A dlycontrol4_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_delay_sample_n12_in sample_n_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[0\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_B edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_307 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[1\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_156 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[2\]
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[3\]
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_17_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[3\]
+ dlycontrol4_in[3] VSS VDD sky130_fd_sc_hd__inv_2
XPHY_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A dlycontrol1_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_delay_sample_p11_in sample_p_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_226 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1 clkgen.clk_dig_out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_270 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_211 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A dlycontrol2_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XPHY_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[3\]
+ dlycontrol3_in[3] VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_225 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_280 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_3.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_6_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_195 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A dlycontrol3_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_259 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_292 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_9_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_A1 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_268 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[4\]
+ dlycontrol1_in[4] VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A dlycontrol4_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_216 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_263 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_226 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VSS VDD sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
.ends

.subckt sky130_fd_sc_hd__dfstp_2 VPWR VGND Q SET_B D CLK VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X15 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X20 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X21 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.21 as=0.12075 ps=1.165 w=0.84 l=0.15
X24 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X25 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X27 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X28 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X29 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt adc_top clk_vcm config_1_in[0] config_1_in[10] config_1_in[11] config_1_in[12]
+ config_1_in[13] config_1_in[14] config_1_in[15] config_1_in[1] config_1_in[2] config_1_in[3]
+ config_1_in[4] config_1_in[5] config_1_in[6] config_1_in[7] config_1_in[8] config_1_in[9]
+ config_2_in[0] config_2_in[10] config_2_in[11] config_2_in[12] config_2_in[13] config_2_in[14]
+ config_2_in[15] config_2_in[1] config_2_in[2] config_2_in[3] config_2_in[4] config_2_in[5]
+ config_2_in[6] config_2_in[7] config_2_in[8] config_2_in[9] conversion_finished_osr_out
+ conversion_finished_out inn_analog inp_analog result_out[0] result_out[10] result_out[11]
+ result_out[12] result_out[13] result_out[14] result_out[15] result_out[1] result_out[2]
+ result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8]
+ result_out[9] rst_n start_conversion_in VDD VSS
X_3155_ VSS VDD net59 _0045_ net71 net40 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3086_ VDD VSS _1342_ _0971_ _0799_ VSS VDD sky130_fd_sc_hd__xor2_1
X_2106_ VDD VSS _1125_ _0068_ core.pdc.col_out\[27\] _0070_ _1102_ _0160_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
X_2037_ VDD VSS _0120_ _0098_ VSS VDD sky130_fd_sc_hd__inv_2
X_2939_ VSS VDD _0830_ _0831_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1534__A net15 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3132__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_93_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2084__B _0113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_83_309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1987__A2 _1053_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2724_ VSS VDD _0620_ _0622_ _0621_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2655_ VSS VDD _0288_ _0560_ _0530_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1606_ VDD VSS _1154_ _1153_ VSS VDD sky130_fd_sc_hd__inv_2
X_2586_ VSS VDD _1300_ _0501_ _0502_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1537_ VSS VDD _1075_ _1084_ _1070_ _1064_ core.ndc.col_out_n\[1\] _1094_ VSS VDD
+ sky130_fd_sc_hd__o221a_2
X_1468_ VSS VDD _1028_ _1030_ _1029_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3138_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0028_ net85 core.cnb.result_out\[6\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3069_ VDD VSS _0955_ _0954_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_88_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2095__A _0065_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1439__A _1002_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[3\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[3\] core.pdc.row_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__3178__CLK net58 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2440_ VSS VDD _1332_ core.pdc.rowon_bottotop_n\[5\] _1342_ VSS VDD sky130_fd_sc_hd__nor2_2
X_2371_ VSS VDD _0384_ core.osr.result_r\[18\] _0387_ VSS VDD sky130_fd_sc_hd__nand2b_1
XFILLER_56_309 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1902__A core.pdc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2082__A1 _1284_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2707_ VSS VDD _0376_ _0605_ _0606_ _0517_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_2638_ VSS VDD core.osr.next_result_w\[7\] _0545_ _0535_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2569_ VSS VDD _1395_ _0483_ _0490_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_59_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2908__A _0799_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_489 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_130_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_31 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2362__B _0241_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_139_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_99_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_99_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_9_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1940_ VSS VDD _1396_ _1395_ _1394_ _1079_ _1085_ VSS VDD sky130_fd_sc_hd__a211o_2
X_1871_ VSS VDD core.ndc.rowoff_out_n\[8\] _1321_ _1352_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2423_ VSS VDD _1356_ _1352_ core.ndc.row_out_n\[4\] VSS VDD sky130_fd_sc_hd__nor2_1
X_2354_ VSS VDD _0371_ _0373_ _0372_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2285_ VSS VDD _0309_ _0311_ _0307_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2447__B core.pdc.rowon_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_301 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk2\[0\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[0\] core.ndc.row_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_100_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2182__B _0220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1802__A1 _1126_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1802__B2 _1296_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_60_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_118_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_118_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_109_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1807__A core.cnb.data_register_r\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_183 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_34_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2267__B core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2070_ VDD VSS core.pdc.col_out_n\[18\] core.pdc.col_out\[18\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1598__S _1077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2972_ VSS VDD _0054_ _0757_ _0863_ _0861_ _1055_ _0688_ VSS VDD sky130_fd_sc_hd__a32o_1
X_1923_ VSS VDD _1362_ core.ndc.rowoff_out_n\[5\] _1384_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1854_ VSS VDD _1340_ _1026_ _1341_ _1300_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1627__A _1032_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1785_ VSS VDD _1124_ _1291_ _1275_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2406_ VDD VSS _0414_ core.osr.is_last_sample _0412_ _0415_ VSS VDD sky130_fd_sc_hd__or3_1
X_2337_ VDD VSS _0358_ _0357_ VSS VDD sky130_fd_sc_hd__inv_2
X_2268_ VSS VDD _0296_ _0294_ _0255_ _0293_ _0295_ VSS VDD sky130_fd_sc_hd__a31o_1
Xgenblk2\[4\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[4\] core.pdc.rowon_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2199_ VSS VDD core.cnb.next_average_sum_w\[3\] _0234_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA_nmat_col_n[8] nmatrix_col_core_n_buffered\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_197 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_136_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_96_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1711__A0 _1242_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input18_A config_2_in[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1570_ VSS VDD _1058_ _1037_ _1122_ VSS VDD sky130_fd_sc_hd__nor2_1
X_3171_ VSS VDD net61 core.osr.next_result_w\[11\] net73 core.osr.result_r\[11\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2122_ VSS VDD _1396_ _0171_ _1188_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_19_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_481 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2053_ VDD VSS _0131_ _0132_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_34_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2955_ VDD VSS _0847_ _0471_ VSS VDD sky130_fd_sc_hd__inv_2
X_1906_ VDD VSS _1376_ _1375_ VSS VDD sky130_fd_sc_hd__inv_2
X_2886_ VSS VDD _0780_ _0777_ _0779_ VSS VDD sky130_fd_sc_hd__or2_1
X_1837_ VSS VDD core.cnb.data_register_r\[10\] _1326_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1768_ VSS VDD _1176_ _1280_ _1279_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1699_ VDD VSS _1232_ _1233_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_85_510 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_122_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2249__A1 core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1820__A _1312_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_101 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_25_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3160__RESET_B net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[8\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[8\] core.pdc.row_out_n\[8\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xoutput42 VDD VSS result_out[13] net42 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput53 VDD VSS result_out[9] net53 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2098__A _0065_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1999__B1 _1259_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2740_ VSS VDD _0206_ _0636_ _0635_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2561__A _0482_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2671_ VSS VDD _0347_ _1002_ _0574_ _0348_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_75_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1622_ VDD VSS _1167_ _1168_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_1553_ VDD VSS core.ndc.col_out_n\[2\] core.ndc.col_out\[2\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2500__S _0220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1484_ VDD VSS _1044_ core.cnb.data_register_r\[5\] VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1624__B _1045_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3154_ VSS VDD net59 _0044_ net71 net39 VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__1640__A _1039_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3085_ VSS VDD _0966_ _0970_ _0969_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2105_ VDD VSS _0160_ _0103_ _1092_ VSS VDD sky130_fd_sc_hd__and2_1
X_2036_ VSS VDD _0118_ _0119_ _1235_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2938_ VSS VDD _0820_ _0829_ _0830_ _0753_ VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__2471__A core.pdc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2869_ VSS VDD _0649_ _0701_ _0763_ _0762_ VSS VDD sky130_fd_sc_hd__nand3_1
Xgenblk1\[3\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[3\] core.pdc.col_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1914__B1 core.ndc.rowon_bottotop_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_42_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2381__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1709__B _1213_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_67_82 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk2\[5\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[5\] core.ndc.row_bottotop_n\[5\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2723_ VDD VSS _0530_ _0356_ _1018_ _0621_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_2654_ VSS VDD _0557_ _0559_ _0558_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1605_ VSS VDD _1105_ _1078_ _1153_ _1135_ VSS VDD sky130_fd_sc_hd__a21oi_2
X_2585_ VSS VDD _0488_ _0501_ _1067_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1635__A core.ndc.col_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1536_ VSS VDD _1091_ _1094_ _1093_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1467_ VSS VDD core.cnb.data_register_r\[11\] _1029_ core.cnb.data_register_r\[10\]
+ VSS VDD sky130_fd_sc_hd__nor2_2
X_3137_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0027_ net79 core.cnb.result_out\[5\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_3068_ VDD VSS _1326_ _0954_ _0799_ VSS VDD sky130_fd_sc_hd__xor2_1
X_2019_ VSS VDD _0107_ _0108_ _1135_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_50_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1545__A _1032_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_92_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2823__B core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[0\].buf_n_coln VDD VSS core.ndc.col_out_n\[0\] nmatrix_col_core_n_buffered\[0\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_2370_ VSS VDD core.osr.next_result_w\[17\] _0386_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_68_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1902__B _1325_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3122__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2706_ VSS VDD _0381_ _0385_ _0605_ _0517_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2637_ VSS VDD core.osr.next_result_w\[9\] _0544_ _0533_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_58_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2568_ VDD VSS _0489_ _0488_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_2499_ VSS VDD _0004_ _0440_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1519_ VDD VSS _1077_ _1041_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_114_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_114_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_56 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_99_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_99_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_405 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1722__B _1102_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1870_ VDD VSS core.ndc.rowoff_out_n\[8\] _1351_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_80_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2422_ VSS VDD _1350_ _1354_ core.ndc.row_out_n\[3\] VSS VDD sky130_fd_sc_hd__nor2_1
X_2353_ VSS VDD _0352_ _0372_ _0370_ VSS VDD sky130_fd_sc_hd__or2b_1
X_2284_ VSS VDD _0310_ _0307_ _0309_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1632__B _1177_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1999_ VSS VDD _1259_ _0090_ _0088_ _1224_ core.pdc.col_out_n\[7\] _0093_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_109_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3185__RESET_B net87 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3168__CLK net66 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_195 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_34_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_59_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_151 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2971_ VSS VDD _0862_ _0790_ _0863_ _0805_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1922_ VSS VDD _1372_ _1369_ _1378_ core.pdc.rowon_out_n\[12\] VSS VDD sky130_fd_sc_hd__a21o_2
X_1853_ VSS VDD _1340_ _1339_ _1303_ VSS VDD sky130_fd_sc_hd__nand2_2
XANTENNA__1796__A1 _1091_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1796__B2 _1296_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1908__A _1377_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1784_ VDD VSS _1289_ _1290_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_115_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[8\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[8\] core.pdc.col_out_n\[8\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2405_ VDD VSS _0414_ _0413_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2458__B core.ndc.rowon_out_n\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_29_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2336_ VSS VDD core.osr.result_r\[12\] _0357_ core.osr.result_r\[13\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2267_ VDD VSS _0295_ _0251_ core.cnb.result_out\[6\] VSS VDD sky130_fd_sc_hd__and2_1
X_2198_ VSS VDD _0234_ _0233_ _0232_ _0209_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA_nmat_col_n[7] nmatrix_col_core_n_buffered\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_136_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1553__A core.ndc.col_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2368__B _0255_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1711__A1 _1202_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_416 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_83_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1778__A1 _1284_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1728__A core.ndc.col_out_n\[16\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1463__A net14 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_126 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3170_ VSS VDD net61 core.osr.next_result_w\[10\] net73 core.osr.result_r\[10\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2121_ VSS VDD _1401_ _0170_ _1096_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2052_ VSS VDD _1227_ _0094_ _0131_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1910__B _1342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_493 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2954_ VSS VDD _0845_ _0846_ _0475_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1905_ VSS VDD _1038_ _1339_ _1375_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2741__B net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2885_ VSS VDD _0778_ _0779_ _0718_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1836_ VDD VSS _1325_ _1324_ VSS VDD sky130_fd_sc_hd__buf_2
X_1767_ VDD VSS _1279_ _1032_ VSS VDD sky130_fd_sc_hd__buf_2
X_1698_ VSS VDD _1227_ _1231_ _1232_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2497__A2 _0220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2319_ VDD VSS _0342_ _0341_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_66_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_85_522 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1820__B _1022_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[5\].buf_n_coln VDD VSS core.ndc.col_out_n\[5\] nmatrix_col_core_n_buffered\[5\]
+ VSS VDD sky130_fd_sc_hd__buf_6
Xoutput43 VDD VSS result_out[14] net43 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2098__B _0115_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1696__A0 _1229_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input30_A config_2_in[6] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1730__B _1213_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1999__A1 _1224_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_31_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2670_ VDD VSS _1008_ _0363_ _0524_ _0573_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_1621_ VSS VDD _1131_ _1166_ _1167_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1552_ VDD VSS _1096_ core.ndc.col_out\[2\] _1091_ _1107_ _1100_ _1102_ VSS VDD sky130_fd_sc_hd__a221o_4
X_1483_ VSS VDD _1042_ _1043_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3153_ VSS VDD net59 _0043_ net71 net53 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_100_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1921__A _1383_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2104_ VDD VSS core.pdc.col_out\[26\] core.pdc.col_out_n\[26\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_3084_ VDD VSS _0918_ _0912_ _1022_ _0969_ VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_47_290 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2035_ VDD VSS _0118_ _0074_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_22_146 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2937_ VSS VDD _0828_ _0809_ _0806_ _0829_ VSS VDD sky130_fd_sc_hd__nor3_1
XANTENNA__2471__B core.pdc.rowon_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2868_ VSS VDD core.cnb.shift_register_r\[12\] _0698_ _0762_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1819_ VSS VDD _1071_ _1312_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2799_ VDD VSS _0694_ _0678_ core.cnb.shift_register_r\[15\] VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_133_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_85_374 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_42_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1725__B _1177_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1669__A0 _1208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_116 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1741__A _1033_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1460__B core.cnb.data_register_r\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[13\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[13\] core.ndc.rowon_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2722_ VSS VDD _0618_ _0619_ _0620_ _0528_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2653_ VSS VDD core.osr.next_result_w\[11\] _0558_ _0533_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2584_ VSS VDD core.cnb.result_out\[7\] _0461_ _0500_ _0029_ VSS VDD sky130_fd_sc_hd__o21a_1
X_1604_ VDD VSS _1152_ _1092_ VSS VDD sky130_fd_sc_hd__buf_2
X_1535_ VDD VSS _1093_ _1092_ VSS VDD sky130_fd_sc_hd__buf_2
X_1466_ VSS VDD core.cnb.data_register_r\[9\] core.cnb.data_register_r\[8\] _1028_
+ VSS VDD sky130_fd_sc_hd__nor2_1
X_3136_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0026_ net78 core.cnb.result_out\[4\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_55_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3067_ VSS VDD _0952_ _0059_ _0953_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2018_ VSS VDD _1390_ _0107_ _1122_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2482__A core.pdc.row_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_A net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2657__A _0983_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1561__A _1114_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1736__A _1124_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1471__A core.ndc.rowoff_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2705_ VSS VDD _0602_ _0046_ _0604_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2636_ VSS VDD _0038_ _0541_ _0540_ _0539_ _0543_ VSS VDD sky130_fd_sc_hd__a31o_1
XANTENNA__1593__A2 _1141_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2567_ VSS VDD _0487_ _0473_ _0488_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2498_ VSS VDD _0440_ core.cnb.shift_register_r\[3\] _0203_ core.cnb.shift_register_r\[2\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_1518_ VDD VSS _1076_ core.cnb.data_register_r\[3\] VSS VDD sky130_fd_sc_hd__buf_2
X_1449_ VDD VSS _1013_ core.osr.sample_count_r\[7\] VSS VDD sky130_fd_sc_hd__inv_2
Xvcm net1 vcm/phi2 vcm/phi1_n vcm/phi1 vcm/phi2_n vcm/vcm VDD vcm/mimtop1 vcm/mimtop2
+ vcm/mimbot1 VSS adc_vcm_generator
XFILLER_55_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3119_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0019_ net84 core.cnb.sampled_avg_control_r\[0\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_82_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_130_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_11 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_99_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1556__A _1039_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_417 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_104_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_80_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2421_ VSS VDD _1331_ _1329_ core.ndc.row_out_n\[2\] _1357_ VSS VDD sky130_fd_sc_hd__a21oi_2
XFILLER_89_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2352_ VSS VDD _0309_ _0351_ _0371_ _0370_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2283_ VSS VDD _0308_ _0300_ _0309_ _0294_ VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_52_358 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_100_49 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1998_ VSS VDD _0092_ _0093_ _1155_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_133_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2619_ VSS VDD _1011_ _0528_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_87_200 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_125_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_125_79 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_461 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2373__C _0240_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2451__B1 _1328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_380 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_108 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3112__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2970_ VSS VDD _0792_ _0862_ _0789_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1921_ VSS VDD core.pdc.rowon_out_n\[11\] _1383_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_98_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_71 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1852_ VDD VSS _1339_ _1338_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1796__A2 _1279_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1783_ VSS VDD _1131_ _1194_ _1289_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2404_ VSS VDD _0410_ _0413_ core.osr.sample_count_r\[5\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2335_ VDD VSS _0356_ core.osr.next_result_w\[12\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2266_ VSS VDD _0292_ _0294_ _0291_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2197_ VSS VDD _0227_ _0233_ core.cnb.average_sum_r\[3\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col_n[6] nmatrix_col_core_n_buffered\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_144 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1834__A _1323_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3135__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_29_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2665__A core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_45_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2120_ VDD VSS core.pdc.col_out_n\[29\] core.pdc.col_out\[29\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_86_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2051_ VSS VDD _1396_ _0130_ _1152_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_47_461 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2953_ VSS VDD _0844_ _0845_ _0834_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1904_ VSS VDD _1374_ _1026_ _1373_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1638__B _1053_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2884_ VSS VDD _0718_ _0720_ _0778_ _0719_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1835_ VSS VDD net14 _1324_ _1308_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1766_ VDD VSS core.ndc.col_out\[23\] core.ndc.col_out_n\[23\] VSS VDD sky130_fd_sc_hd__inv_2
X_1697_ VDD VSS _1231_ _1230_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_106_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2318_ VSS VDD core.osr.result_r\[11\] _0341_ core.cnb.result_out\[11\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2249_ VSS VDD _0278_ core.cnb.result_out\[4\] _0279_ _0271_ VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_82_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_89 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1829__A _1022_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[0\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[0\] core.pdc.rowon_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xoutput44 VDD VSS result_out[15] net44 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1696__A1 _1161_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input23_A config_2_in[14] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_515 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_56_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1739__A core.ndc.col_out_n\[18\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1620_ VDD VSS _1166_ _1165_ VSS VDD sky130_fd_sc_hd__inv_2
X_1551_ VDD VSS _1107_ _1106_ _1092_ VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__1474__A _1033_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1482_ VDD VSS _1042_ _1041_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_97_92 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_309 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3152_ VSS VDD net57 _0042_ net69 net52 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2103_ VDD VSS _1152_ _0146_ core.pdc.col_out\[26\] _0118_ _1102_ _0159_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
X_3083_ VSS VDD _0967_ _0968_ _0060_ _0758_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_2034_ VDD VSS _0116_ _0117_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_50_423 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_445 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_489 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2936_ VSS VDD _0825_ _0726_ _0828_ _0827_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2867_ VSS VDD _0471_ _0761_ _0760_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1818_ VDD VSS _1310_ _1311_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_2798_ VSS VDD _0640_ _0660_ _0693_ _0454_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_117_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1749_ VSS VDD _1212_ _1269_ _1177_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_133_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_26_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_13_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_512 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1669__A1 _1197_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[14\].buf_p_rowonn_A core.pdc.rowon_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3014__A _1312_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1469__A net14 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2721_ VSS VDD core.osr.next_result_w\[18\] _0619_ _0533_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2652_ VDD VSS core.osr.next_result_w\[9\] _0535_ _0556_ _0557_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_1603_ VDD VSS core.ndc.col_out_n\[5\] core.ndc.col_out\[5\] VSS VDD sky130_fd_sc_hd__inv_2
X_2583_ VDD VSS _0489_ _1067_ _0500_ _0498_ _1117_ _0439_ VSS VDD sky130_fd_sc_hd__a221o_1
X_1534_ VSS VDD net15 _1092_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1465_ VSS VDD core.ndc.rowoff_out_n\[0\] _1025_ _1027_ VSS VDD sky130_fd_sc_hd__nand2_2
X_3204_ VSS VDD net65 core.osr.is_last_sample net84 core.osr.data_valid_r VSS VDD
+ sky130_fd_sc_hd__dfrtp_1
X_3135_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0025_ net78 core.cnb.result_out\[3\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3066_ VSS VDD _0758_ _0953_ _1303_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2017_ VSS VDD _0106_ _1133_ _1390_ _1137_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__2482__B core.pdc.rowon_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2919_ VSS VDD _0810_ _0730_ _0811_ _0731_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_128_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_128_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_fanout73_A net83 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1561__B _1037_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_68_117 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1471__B core.ndc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1927__A core.ndc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2704_ VDD VSS _0604_ _0603_ VSS VDD sky130_fd_sc_hd__inv_2
X_2635_ VDD VSS _0394_ core.cnb.result_out\[0\] _0542_ _0543_ net48 VSS VDD sky130_fd_sc_hd__a22o_1
X_2566_ VDD VSS core.cnb.data_register_r\[0\] _0482_ _1076_ core.cnb.data_register_r\[1\]
+ _0487_ VSS VDD sky130_fd_sc_hd__or4_1
X_1517_ VDD VSS _1075_ _1074_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_59_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2497_ VSS VDD _0220_ _0439_ _0003_ _0437_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__2477__B core.pdc.row_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1448_ VSS VDD _1011_ _1012_ _0985_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3118_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0018_ net86 core.cnb.shift_register_r\[16\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_130_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3049_ VSS VDD _0882_ _0868_ _0937_ _0906_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_90_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_139_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_rowoff_n[1] core.ndc.rowoff_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout90 VSS VDD net92 net90 VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1747__A _1187_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1466__B core.cnb.data_register_r\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2420_ VSS VDD _1344_ _1359_ core.ndc.row_out_n\[1\] VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1980__B1 _1259_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3191__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2351_ VSS VDD _0370_ core.osr.result_r\[15\] core.osr.result_r\[14\] _0358_ VSS
+ VDD sky130_fd_sc_hd__and3_1
X_2282_ VSS VDD _0290_ _0297_ _0298_ _0308_ VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_92_440 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_92_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1997_ VDD VSS _0092_ _0091_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_133_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2618_ VSS VDD _0519_ core.osr.next_result_w\[3\] _0527_ core.osr.next_result_w\[7\]
+ _0526_ _0524_ VSS VDD sky130_fd_sc_hd__o221ai_1
X_2549_ VSS VDD _0472_ _0438_ _0473_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_87_212 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_56 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_115_91 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1920_ VSS VDD _1383_ _1382_ _1373_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_91_83 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2861__A _0691_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1851_ VSS VDD _1338_ _1326_ core.cnb.data_register_r\[11\] VSS VDD sky130_fd_sc_hd__nand2_2
X_1782_ VDD VSS core.ndc.col_out_n\[26\] core.ndc.col_out\[26\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_115_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2403_ VSS VDD core.osr.sample_count_r\[5\] _0410_ _0412_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2334_ VSS VDD _0355_ _0354_ _0356_ _0241_ VSS VDD sky130_fd_sc_hd__nand3_2
X_2265_ VSS VDD _0293_ _0291_ _0292_ VSS VDD sky130_fd_sc_hd__or2_1
X_2196_ VSS VDD _0228_ _0232_ _0231_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_52_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_111_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_nmat_col_n[5] nmatrix_col_core_n_buffered\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_20_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_genblk1\[7\].buf_n_coln_A core.ndc.col_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2011__A _0101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1760__A _1131_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2050_ VDD VSS core.pdc.col_out_n\[14\] core.pdc.col_out\[14\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA_genblk2\[12\].buf_p_rown_A core.pdc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2952_ VSS VDD _0842_ _0844_ _0843_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1903_ VSS VDD _1342_ _1327_ _1373_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2883_ VDD VSS _0777_ _0776_ VSS VDD sky130_fd_sc_hd__inv_2
X_1834_ VDD VSS core.pdc.row_out_n\[3\] _1323_ VSS VDD sky130_fd_sc_hd__inv_2
X_1765_ VSS VDD core.ndc.col_out_n\[23\] _1278_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2530__S net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1696_ VSS VDD _1230_ _1161_ _1041_ _1229_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2317_ VSS VDD core.osr.result_r\[11\] core.cnb.result_out\[11\] _0340_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2248_ VDD VSS _0277_ _0276_ _0252_ _0278_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__1670__A _1033_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2179_ VDD VSS _0218_ core.cnb.average_sum_r\[0\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_25_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__3102__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1564__B _1117_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput45 VDD VSS result_out[1] net45 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2676__A _0395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1580__A core.ndc.col_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input16_A config_1_in[8] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_56_281 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1550_ VSS VDD _1106_ _1105_ _1104_ _1103_ _1088_ VSS VDD sky130_fd_sc_hd__a31o_1
XANTENNA_pmat_col[31] core.pdc.col_out\[31\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1481_ VSS VDD _1041_ core.ndc.rowon_out_n\[0\] _1040_ VSS VDD sky130_fd_sc_hd__nand2_2
X_3151_ VSS VDD net57 _0041_ net71 net51 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2102_ VDD VSS _0159_ _0158_ VSS VDD sky130_fd_sc_hd__inv_2
X_3082_ VSS VDD _0758_ _0968_ _1326_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2033_ VSS VDD _1033_ _0115_ _0116_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__3125__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2935_ VSS VDD _0826_ _0731_ _0827_ _0725_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2866_ VDD VSS _0760_ _0759_ VSS VDD sky130_fd_sc_hd__inv_2
X_1817_ VSS VDD _1309_ _1038_ _1310_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1665__A core.ndc.col_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2797_ VSS VDD _0471_ _0692_ _0686_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1748_ VSS VDD _1221_ _1268_ _1173_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_89_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_117_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1679_ VDD VSS _1217_ _1198_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_input8_A config_1_in[15] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2496__A _0438_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_13_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1850__A2 _1312_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1575__A _1053_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_101_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xgenblk2\[11\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[11\] core.pdc.row_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_49_524 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2720_ VDD VSS _0568_ core.osr.next_result_w\[14\] _0617_ _0618_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_80_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2651_ VDD VSS _1001_ core.osr.next_result_w\[7\] _0530_ _0556_ VSS VDD sky130_fd_sc_hd__a21o_1
X_1602_ VSS VDD _1151_ core.ndc.col_out\[5\] VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2582_ VDD VSS core.cnb.result_out\[6\] _0439_ _0028_ _0497_ _1104_ _0499_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
X_1533_ VSS VDD _1078_ _1090_ _1086_ _1091_ VSS VDD sky130_fd_sc_hd__mux2_2
X_1464_ VSS VDD _1026_ _1027_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3203_ VSS VDD net65 _0064_ net78 core.osr.osr_mode_r\[2\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3134_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0024_ net78 core.cnb.result_out\[2\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_55_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3065_ VSS VDD _0950_ _0781_ _0952_ _0951_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2016_ VDD VSS core.pdc.col_out_n\[9\] core.pdc.col_out\[9\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_50_221 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_107 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2918_ VSS VDD _0638_ _0706_ _0810_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2849_ VSS VDD _0744_ _0645_ _0644_ _0654_ _0650_ VSS VDD sky130_fd_sc_hd__and4_1
XANTENNA_nmat_sample_n _0001_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout66_A net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_68_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_73_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2703_ VDD VSS core.osr.next_result_w\[8\] net41 _1020_ _0603_ _0562_ VSS VDD sky130_fd_sc_hd__a22o_1
X_2634_ VSS VDD _0983_ _0542_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2565_ VSS VDD _0024_ _0486_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1516_ VSS VDD _1073_ _1074_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2496_ VSS VDD _0438_ _0439_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1447_ VDD VSS _1011_ _1009_ VSS VDD sky130_fd_sc_hd__inv_2
X_3117_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0017_ net93 core.cnb.shift_register_r\[15\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__2774__A _0637_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_368 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3048_ VSS VDD _0909_ _0922_ _0936_ _0935_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_64_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_139_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_114 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_nmat_rowoff_n[0] core.ndc.rowoff_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xfanout91 VDD VSS net91 net92 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout80 VDD VSS net80 net81 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2221__A2 _0240_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1747__B _1152_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1980__A1 _1224_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2859__A core.cnb.pswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2350_ VSS VDD _0366_ _0369_ _0368_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2281_ _0307_ _0305_ _0306_ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA__1799__B2 _1296_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1799__A1 _1121_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1996_ VSS VDD _1045_ _1169_ _0091_ _1409_ VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_133_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2617_ VSS VDD _0288_ _0526_ _1002_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1673__A _1092_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2548_ VDD VSS _0471_ _0472_ VSS VDD sky130_fd_sc_hd__buf_6
Xgenblk1\[12\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[12\] core.pdc.col_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2479_ VSS VDD core.pdc.rowon_out_n\[12\] core.pdc.rowoff_out_n\[12\] core.pdc.row_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_18_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1848__A _1335_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_131_91 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2861__B _0208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1850_ VSS VDD _1337_ _1309_ _1312_ _1332_ _1336_ VSS VDD sky130_fd_sc_hd__a31o_1
X_1781_ VSS VDD _1035_ _1143_ _1220_ _1259_ core.ndc.col_out_n\[26\] _1288_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
X_2402_ VDD VSS _0411_ core.osr.next_sample_count_w\[4\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2333_ VSS VDD _0353_ _0355_ core.osr.result_r\[12\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2902__B1 _1076_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2101__B _1072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2264_ VSS VDD _0286_ _0292_ _0282_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2195_ VDD VSS _0231_ core.cnb.average_sum_r\[3\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_52_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[4] nmatrix_col_core_n_buffered\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_179 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1668__A _1206_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1979_ VSS VDD _0077_ _0078_ _1155_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_121_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[6\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[6\] core.ndc.rowon_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2011__B _1275_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_11 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_43_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_43_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__3181__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1578__A _1126_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1760__B _1243_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2951_ VSS VDD _0753_ _0843_ VSS VDD sky130_fd_sc_hd__clkinvlp_2
X_1902_ VSS VDD core.pdc.rowoff_out_n\[5\] core.pdc.rowon_out_n\[4\] _1325_ VSS VDD
+ sky130_fd_sc_hd__nand2_1
X_2882_ VSS VDD _0774_ _0776_ _0775_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1833_ VSS VDD _1322_ core.pdc.rowoff_out_n\[8\] _1323_ _1321_ VSS VDD sky130_fd_sc_hd__o21ai_2
X_1764_ VSS VDD _1278_ _1277_ _1276_ _1274_ VSS VDD sky130_fd_sc_hd__and3_1
X_1695_ VSS VDD _1136_ _1229_ _1228_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2316_ VSS VDD _0338_ _0339_ _0328_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2247_ VSS VDD _0275_ _0277_ _0274_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_122_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2103__A1 _1152_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2103__B2 _1102_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2178_ VSS VDD core.cnb.next_average_counter_w\[4\] _0217_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_53_466 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_68 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_31_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1917__A1 core.ndc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput46 VDD VSS result_out[2] net46 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_56_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_56_293 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1605__B1 _1135_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2030__B1 _1259_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[13\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[13\] core.ndc.row_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1480_ VSS VDD _1040_ _1038_ _1039_ VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_98_116 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3150_ VSS VDD net57 _0040_ net69 net50 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3081_ VSS VDD _0965_ _0691_ _0967_ _0966_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2101_ VSS VDD _0077_ _0158_ _1072_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2032_ VSS VDD _1389_ _1201_ _1199_ _0115_ VSS VDD sky130_fd_sc_hd__mux2_2
X_2934_ VSS VDD _0826_ _0762_ _0645_ _0722_ VSS VDD sky130_fd_sc_hd__and3_1
X_2865_ VSS VDD _0677_ _0713_ _0759_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1816_ VDD VSS _1309_ _1308_ VSS VDD sky130_fd_sc_hd__buf_2
X_2796_ VSS VDD core.cnb.data_register_r\[0\] _0690_ _0687_ _0210_ _0050_ _0691_ VSS
+ VDD sky130_fd_sc_hd__o221a_1
XANTENNA__2021__B1 _1064_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1747_ VSS VDD _1187_ _1267_ _1152_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1678_ VDD VSS core.ndc.col_out\[10\] core.ndc.col_out_n\[10\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2012__A0 _1186_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2618__A2 core.osr.next_result_w\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2079__B1 _1125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2650_ VDD VSS _0554_ _0553_ _0555_ _0040_ VSS VDD sky130_fd_sc_hd__a21o_1
X_1601_ VSS VDD _1144_ _1150_ _1140_ _1151_ VSS VDD sky130_fd_sc_hd__or3b_1
X_2581_ VSS VDD _0439_ _0498_ _0499_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1532_ VSS VDD _1036_ _1089_ _1090_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1463_ VDD VSS _1026_ net14 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_3202_ VSS VDD net64 _0063_ net78 core.osr.osr_mode_r\[1\] VSS VDD sky130_fd_sc_hd__dfrtp_1
Xgenblk1\[17\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[17\] core.pdc.col_out_n\[17\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_55_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3133_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0023_ net84 core.cnb.result_out\[1\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_94_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3064_ VSS VDD _0942_ _0902_ _0951_ _0948_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2015_ VDD VSS core.pdc.col_out_n\[9\] _0105_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_380 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2917_ VSS VDD _0454_ _0808_ _0809_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_12_59 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2848_ VSS VDD _0738_ _0742_ _0743_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2779_ VSS VDD _0672_ _0675_ _0674_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__3188__RESET_B net87 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_517 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout59_A net61 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1586__A _1135_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_78_63 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_78_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3115__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_76_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2702_ VSS VDD _0599_ _0602_ _0601_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2633_ VSS VDD _0541_ _0537_ core.osr.next_result_w\[2\] VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_57_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2564_ VSS VDD _0486_ core.cnb.result_out\[2\] _0480_ _0485_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1515_ VDD VSS _1073_ _1072_ VSS VDD sky130_fd_sc_hd__inv_2
X_2495_ VSS VDD _0438_ _0208_ core.cnb.shift_register_r\[2\] VSS VDD sky130_fd_sc_hd__nand2_2
X_1446_ VSS VDD _1009_ _1010_ core.osr.sample_count_r\[2\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_2_3__f_clk_dig_dummy_A clknet_0_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_130 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_325 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3116_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0016_ net93 core.cnb.shift_register_r\[14\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_82_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3047_ VSS VDD _0934_ _0935_ _0906_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_130_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__3097__S _0241_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[14\].buf_n_coln VDD VSS core.ndc.col_out_n\[14\] nmatrix_col_core_n_buffered\[14\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__2949__B _0482_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3138__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_58_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_314 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_73_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[14\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[14\] core.pdc.rowon_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_54_380 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_120_60 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_80_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xfanout92 VDD VSS net92 net94 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout70 VSS VDD net83 net70 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout81 VDD VSS net81 net82 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_127_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2205__A core.cnb.result_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1763__B _1188_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2280_ VSS VDD core.osr.result_r\[8\] _0306_ core.cnb.result_out\[8\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_29_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_453 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_339 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1995_ VDD VSS _0090_ _0089_ VSS VDD sky130_fd_sc_hd__inv_2
X_2616_ VDD VSS _0523_ net46 _0395_ _0036_ _0525_ VSS VDD sky130_fd_sc_hd__a22o_1
XANTENNA__1954__A _1272_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2547_ VDD VSS _0470_ _0471_ VSS VDD sky130_fd_sc_hd__buf_6
X_2478_ VSS VDD core.pdc.row_out_n\[11\] core.pdc.rowoff_out_n\[11\] core.pdc.rowon_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1429_ VSS VDD core.osr.osr_mode_r\[2\] _0989_ _0993_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_18_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_361 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2025__A _0101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_109_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_93_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_131_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xnmat_sample_buf VSS VDD nmat_sample_switch_buffered net55 VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_91_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1780_ VSS VDD _1149_ _1288_ _1284_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1774__A _1095_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2401_ VDD VSS _0410_ core.osr.is_last_sample _0409_ _0411_ VSS VDD sky130_fd_sc_hd__or3_1
X_2332_ VSS VDD _0354_ core.osr.result_r\[12\] _0353_ VSS VDD sky130_fd_sc_hd__or2_1
X_2263_ VDD VSS _0291_ _0289_ _0290_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_84_228 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2194_ VSS VDD core.cnb.next_average_sum_w\[2\] _0230_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_92_261 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col_n[3] nmatrix_col_core_n_buffered\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1978_ VSS VDD _0077_ _1146_ _1400_ _1147_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_121_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col[19] core.ndc.col_out\[19\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_409 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_29_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_144 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_90_209 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_83_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1859__A _1325_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1578__B _1129_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_101_84 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1594__A _1074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_120_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1533__S _1078_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2950_ VSS VDD _0832_ _0842_ _0833_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1488__B _1047_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1901_ VSS VDD core.pdc.rowoff_out_n\[5\] _1372_ _1309_ VSS VDD sky130_fd_sc_hd__nand2_2
X_2881_ VSS VDD _0771_ _0772_ _0775_ _0482_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1832_ VDD VSS _1308_ _1304_ _1038_ _1300_ _1322_ VSS VDD sky130_fd_sc_hd__or4_1
X_1763_ VSS VDD _1180_ _1277_ _1188_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1694_ VDD VSS _1228_ _1105_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_106_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2315_ VSS VDD _0326_ _0338_ _0330_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2246_ VSS VDD _0276_ _0274_ _0275_ VSS VDD sky130_fd_sc_hd__or2_1
X_2177_ VSS VDD _0217_ _0216_ _0215_ _0210_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_25_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_1__leaf_clk_dig_dummy
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xgenblk1\[24\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[24\] core.pdc.col_out_n\[24\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xoutput47 VDD VSS result_out[3] net47 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput36 VDD VSS conversion_finished_osr_out net36 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2957__B core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1550__B1 _1088_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_56_99 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_56_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1589__A _1138_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk1\[3\].buf_n_coln_A core.ndc.col_out_n\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1605__A1 _1078_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2030__A1 _1074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3080_ VSS VDD _0964_ _0966_ _0955_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2100_ VDD VSS core.pdc.col_out_n\[25\] core.pdc.col_out\[25\] VSS VDD sky130_fd_sc_hd__inv_2
X_2031_ VDD VSS core.pdc.col_out_n\[12\] core.pdc.col_out\[12\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_22_106 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2933_ VSS VDD _0821_ _0824_ _0825_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_87_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2864_ VSS VDD _0051_ _0757_ _0755_ _0721_ core.cnb.data_register_r\[1\] _0758_ VSS
+ VDD sky130_fd_sc_hd__a32o_1
X_1815_ VSS VDD core.cnb.data_register_r\[11\] _1308_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2795_ VSS VDD _0460_ _0691_ _0670_ VSS VDD sky130_fd_sc_hd__nor2_2
XANTENNA__1946__B _1155_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1746_ VDD VSS core.ndc.col_out\[19\] core.ndc.col_out_n\[19\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2021__A1 _1224_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2123__A _1039_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1677_ VSS VDD _1216_ core.ndc.col_out_n\[10\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__3171__CLK net61 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[19\].buf_n_coln VDD VSS core.ndc.col_out_n\[19\] nmatrix_col_core_n_buffered\[19\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__1681__B _1173_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_312 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2229_ VSS VDD _0259_ _0261_ _0258_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_26_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2796__C1 _0691_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2012__A1 _1197_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2033__A _1033_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_107_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_67_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_input21_A config_2_in[12] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2079__A1 _1102_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_91_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2208__A _0241_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[21\].buf_n_coln VDD VSS core.ndc.col_out_n\[21\] nmatrix_col_core_n_buffered\[21\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_83_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1600_ VSS VDD _1149_ _1150_ _1032_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2580_ VSS VDD _0489_ _0498_ _1160_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1531_ VDD VSS _1089_ _1088_ VSS VDD sky130_fd_sc_hd__inv_2
X_1462_ VSS VDD _1024_ _1025_ core.cnb.data_register_r\[11\] VSS VDD sky130_fd_sc_hd__nand2_1
X_3201_ VSS VDD net65 _0062_ net78 core.osr.osr_mode_r\[0\] VSS VDD sky130_fd_sc_hd__dfrtp_2
X_3132_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0022_ net84 core.cnb.result_out\[0\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_3063_ VSS VDD _0944_ _0950_ _0949_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2014_ VSS VDD _0105_ _0104_ _0102_ _0100_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_90_392 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2916_ VSS VDD _0807_ _0808_ _0725_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2847_ VSS VDD _0742_ _0649_ _0724_ _0741_ VSS VDD sky130_fd_sc_hd__and3_1
X_2778_ VSS VDD _0674_ _0640_ _0652_ _0673_ VSS VDD sky130_fd_sc_hd__nand3b_1
XANTENNA__1692__A core.ndc.col_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1729_ VSS VDD _1255_ _1074_ _1243_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_37_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_507 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1992__B1 _1082_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_78_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_78_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_76_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_134 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2880__B core.cnb.pswitch_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2701_ VDD VSS _0601_ _0600_ VSS VDD sky130_fd_sc_hd__inv_2
X_2632_ VSS VDD _1019_ _0540_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2563_ VSS VDD _0483_ _0485_ _0484_ VSS VDD sky130_fd_sc_hd__or2b_1
X_1514_ VSS VDD _1071_ _1072_ net15 VSS VDD sky130_fd_sc_hd__nor2_2
X_2494_ VDD VSS _0437_ core.cnb.is_holding_result_w VSS VDD sky130_fd_sc_hd__inv_2
X_1445_ VSS VDD _1008_ _1009_ core.osr.osr_mode_r\[1\] VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_67_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3115_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0015_ net93 core.cnb.shift_register_r\[13\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_55_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3046_ VSS VDD _0928_ _0933_ _0934_ _0870_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_82_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout71_A net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout60 VSS VDD net60 net61 VSS VDD sky130_fd_sc_hd__clkbuf_1
Xfanout71 VSS VDD net73 net71 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout82 VDD VSS net82 net83 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_127_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1965__B1 _1125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout93 VDD VSS net93 net94 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_127_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_92_465 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1994_ VSS VDD _1394_ _1242_ _1202_ _0089_ VSS VDD sky130_fd_sc_hd__mux2_2
XANTENNA__2115__B _1096_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[29\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[29\] core.pdc.col_out_n\[29\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2615_ VSS VDD _0525_ _0524_ core.osr.next_result_w\[6\] VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__2131__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2546_ VDD VSS _0469_ _0468_ _0470_ _0203_ VSS VDD sky130_fd_sc_hd__a21boi_2
XFILLER_125_28 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2477_ VSS VDD core.pdc.rowon_out_n\[10\] core.pdc.rowoff_out_n\[10\] core.pdc.row_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1428_ VDD VSS _0992_ _0991_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_18_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3029_ VDD VSS _0916_ _0830_ _0856_ _0917_ VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_51_373 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__3105__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2025__B _1093_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_35 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1947__B1 _1259_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_124_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_59_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xgenblk1\[31\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[31\] core.pdc.col_out_n\[31\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_61_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[1\].buf_n_rown_A core.ndc.row_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2400_ VSS VDD _0999_ _0406_ _0410_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2331_ VSS VDD _0353_ _0351_ _0309_ _0352_ VSS VDD sky130_fd_sc_hd__a21bo_1
X_2262_ VSS VDD core.cnb.result_out\[6\] _0290_ core.osr.result_r\[6\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2193_ VSS VDD _0230_ _0229_ _0228_ _0209_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA_nmat_col_n[2] nmatrix_col_core_n_buffered\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[0\].buf_p_rowonn_A core.pdc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3128__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1977_ VDD VSS _0076_ _0075_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1684__B _1177_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[1\].buf_n_rowonn_A core.ndc.rowon_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col[18] core.ndc.col_out\[18\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2529_ VSS VDD _0018_ _0456_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_29_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_56_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_45_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_43_148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_101_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_181 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[26\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[26\] core.ndc.col_out_n\[26\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_101_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_64 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1769__B _1213_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1900_ VSS VDD _1023_ _1372_ _1022_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2880_ VSS VDD _0773_ _0774_ core.cnb.pswitch_out\[2\] VSS VDD sky130_fd_sc_hd__nand2_1
X_1831_ VSS VDD _1321_ _1318_ core.pdc.rowoff_out_n\[8\] _1311_ core.pdc.row_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__o22a_1
XANTENNA__1785__A _1124_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1762_ VSS VDD _1187_ _1276_ _1275_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1693_ VDD VSS _1227_ _1073_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_103_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_106_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2314_ VDD VSS _0337_ core.osr.next_result_w\[10\] VSS VDD sky130_fd_sc_hd__buf_6
X_2245_ VSS VDD _0267_ _0275_ _0265_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2176_ VSS VDD _0214_ _0216_ core.cnb.average_counter_r\[4\] VSS VDD sky130_fd_sc_hd__nand2_1
Xoutput48 VDD VSS result_out[4] net48 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput37 VDD VSS conversion_finished_out net65 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA_genblk1\[18\].buf_n_coln_A core.ndc.col_out_n\[18\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_398 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1605__A2 _1105_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[2\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[2\] core.ndc.rowon_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA_pmat_col[4] core.pdc.col_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2030__A2 _0113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2030_ VSS VDD _1259_ _0088_ _0113_ _1074_ core.pdc.col_out_n\[12\] _0114_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2932_ VSS VDD _0737_ _0813_ _0824_ _0823_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_94_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2863_ VSS VDD _0688_ _0758_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1814_ VSS VDD _1300_ _1306_ _1307_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2794_ VDD VSS _0690_ _0689_ _0686_ VSS VDD sky130_fd_sc_hd__and2_1
X_1745_ VSS VDD _1266_ core.ndc.col_out_n\[19\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_7_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1676_ VSS VDD _1216_ _1215_ _1214_ _1211_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_85_302 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2228_ VSS VDD _0260_ _0258_ _0259_ VSS VDD sky130_fd_sc_hd__or2_1
X_2159_ VSS VDD _0203_ _0189_ _0202_ VSS VDD sky130_fd_sc_hd__nand2_2
XANTENNA__2796__B1 core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2033__B _0115_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_analog_in ANTENNA_pmat_analog_in/DIODE VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xpmat_95 net95 pmat_95/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_107_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_305 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input14_A config_1_in[6] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1530_ VSS VDD _1088_ _1085_ _1087_ VSS VDD sky130_fd_sc_hd__nor2_4
X_1461_ VSS VDD _1022_ _1023_ _1024_ VSS VDD sky130_fd_sc_hd__nor2_1
X_3200_ VSS VDD net64 core.osr.next_sample_count_w\[8\] net77 core.osr.sample_count_r\[8\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3131_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[4\] net91
+ core.cnb.average_sum_r\[4\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA_genblk2\[5\].buf_p_rowonn_A core.pdc.rowon_bottotop_n\[5\] VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[19] nmatrix_col_core_n_buffered\[19\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3062_ VDD VSS _0949_ _0948_ VSS VDD sky130_fd_sc_hd__inv_2
X_2013_ VSS VDD _0103_ _0104_ _1101_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_76_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2915_ VSS VDD _0807_ _0694_ _0644_ _0722_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_12_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2846_ VSS VDD _0646_ _0634_ _0740_ _0741_ VSS VDD sky130_fd_sc_hd__nor3_1
X_2777_ VSS VDD _0653_ _0673_ core.cnb.shift_register_r\[11\] VSS VDD sky130_fd_sc_hd__nand2_1
X_1728_ VDD VSS core.ndc.col_out\[16\] core.ndc.col_out_n\[16\] VSS VDD sky130_fd_sc_hd__inv_2
X_1659_ VSS VDD _1059_ _1052_ _1201_ _1200_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA_input6_A config_1_in[13] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_37_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_67_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_24 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_53_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1992__A1 _1114_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_136 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_94_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_91_146 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_73_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2700_ VSS VDD core.osr.next_result_w\[10\] _1019_ _0600_ _1011_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1793__A core.ndc.col_out\[28\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2631_ VSS VDD _0534_ _0536_ _0539_ _0538_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2562_ VSS VDD _0478_ _0484_ _0482_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1513_ VDD VSS _1071_ core.cnb.data_register_r\[8\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_4_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2493_ VSS VDD _0220_ _0434_ _0002_ core.cnb.enable_loop_out VSS VDD sky130_fd_sc_hd__o21ai_1
X_1444_ VDD VSS _0993_ _1008_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_3114_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0014_ net93 core.cnb.shift_register_r\[12\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_3045_ VSS VDD _0931_ _1114_ _0933_ _0932_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_64_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2829_ VSS VDD _0642_ _0724_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout64_A net66 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_45 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3184__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_393 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xfanout61 VSS VDD net67 net61 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout72 VDD VSS net72 net73 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout83 VSS VDD net34 net83 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout94 VDD VSS net94 net34 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1965__A1 _1121_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1965__B2 _1413_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_92_477 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1993_ VDD VSS _0088_ _0087_ VSS VDD sky130_fd_sc_hd__inv_2
X_2614_ VSS VDD _0994_ _0524_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2545_ VSS VDD _0469_ _0222_ _0207_ VSS VDD sky130_fd_sc_hd__or2_1
X_2476_ VSS VDD core.pdc.row_out_n\[9\] core.pdc.rowoff_out_n\[9\] core.pdc.rowon_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1427_ VSS VDD _0991_ core.osr.osr_mode_r\[2\] _0990_ _0989_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_83_400 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_83_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3028_ VSS VDD _0916_ _0818_ _0751_ _0910_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_83_477 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1698__A _1227_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1947__A1 _1224_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_47 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk2\[4\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[4\] core.pdc.row_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_93_219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk2\[10\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[10\] core.pdc.rowon_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2330_ VSS VDD _0352_ _0350_ _0342_ _0329_ _0343_ _0324_ VSS VDD sky130_fd_sc_hd__a221oi_1
X_2261_ VSS VDD _0289_ core.cnb.result_out\[6\] core.osr.result_r\[6\] VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_34_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2192_ VSS VDD _0223_ _0229_ _0226_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_37_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col_n[1] nmatrix_col_core_n_buffered\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_296 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1976_ VSS VDD _0075_ _1208_ _1394_ _1197_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__2142__A core.cnb.sampled_avg_control_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_107 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col[17] core.ndc.col_out\[17\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2528_ VSS VDD _0456_ net54 _0219_ _0454_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2459_ VSS VDD core.ndc.rowon_out_n\[4\] core.ndc.rowoff_out_n\[4\] core.ndc.row_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2106__B2 _1102_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2106__A1 _1125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_56_477 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_61_24 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_101_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2036__B _1235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_193 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_61_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2052__A _1227_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_50 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_124 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_34_116 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1830_ VDD VSS _1321_ _1320_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_89_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1785__B _1275_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2584__A1 core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1761_ VDD VSS _1275_ _1072_ VSS VDD sky130_fd_sc_hd__buf_2
X_1692_ VDD VSS core.ndc.col_out\[12\] core.ndc.col_out_n\[12\] VSS VDD sky130_fd_sc_hd__inv_2
Xgenblk2\[1\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[1\] core.ndc.row_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2313_ VDD VSS _0337_ _0334_ _0336_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_25_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2244_ VDD VSS _0274_ _0272_ _0273_ VSS VDD sky130_fd_sc_hd__and2_1
X_2175_ VSS VDD _0215_ core.cnb.average_counter_r\[4\] _0214_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA_cgen_dlycontrol4_in[5] net8 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2024__B1 _1208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2575__A1 core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1959_ VDD VSS _1411_ _1410_ VSS VDD sky130_fd_sc_hd__inv_2
Xoutput49 VDD VSS result_out[5] net49 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput38 VDD VSS result_out[0] net38 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2600__A _1328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_355 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1550__A2 _1104_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_16_116 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2047__A _1413_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_col[3] core.pdc.col_out\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3118__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2931_ VSS VDD _0822_ _0730_ _0823_ _0731_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_30_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2862_ VDD VSS _0757_ _0756_ VSS VDD sky130_fd_sc_hd__inv_2
X_1813_ VSS VDD _1302_ _1306_ _1305_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2793_ VDD VSS _0688_ _0689_ VSS VDD sky130_fd_sc_hd__clkinv_4
X_1744_ VSS VDD _1266_ _1265_ _1264_ _1262_ VSS VDD sky130_fd_sc_hd__and3_1
Xgenblk2\[7\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[7\] core.pdc.rowon_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1675_ VSS VDD _1138_ _1215_ _1177_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2227_ VSS VDD _0249_ _0259_ _0247_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2158_ VSS VDD _0200_ _0202_ _0201_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2089_ VDD VSS _0151_ _0152_ VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__2796__A1 _0210_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_91_317 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_83_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_328 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_60 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1460_ VSS VDD core.cnb.data_register_r\[9\] _1023_ core.cnb.data_register_r\[8\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_79_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3130_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[3\] net91
+ core.cnb.average_sum_r\[3\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_94_100 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[18] nmatrix_col_core_n_buffered\[18\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3061_ VSS VDD _0946_ _0948_ _0947_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2012_ VSS VDD _0103_ _1197_ _1394_ _1186_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2914_ VSS VDD _0806_ _0454_ _0730_ _0725_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__2134__B core.cnb.sampled_avg_control_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2845_ VSS VDD _0653_ _0740_ _0739_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_12_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_128_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2776_ VSS VDD _0669_ _0660_ _0672_ _0671_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1727_ VDD VSS core.ndc.col_out_n\[16\] _1254_ VSS VDD sky130_fd_sc_hd__buf_2
X_1658_ VDD VSS _1200_ _1055_ VSS VDD sky130_fd_sc_hd__inv_2
X_1589_ VDD VSS _1139_ _1138_ VSS VDD sky130_fd_sc_hd__inv_2
Xgenblk2\[9\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[9\] core.pdc.row_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_85_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_37_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_36 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_139_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2325__A core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_158 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2630_ VSS VDD _0519_ _0279_ _0537_ _0538_ VSS VDD sky130_fd_sc_hd__o21a_1
XANTENNA__3066__A _0758_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2561_ VSS VDD _0482_ _0478_ _0483_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2492_ VSS VDD _2492_/X _0436_ VSS VDD sky130_fd_sc_hd__buf_1
X_1512_ VSS VDD _1070_ _1069_ _1054_ _1067_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1443_ VDD VSS _0999_ _0994_ core.osr.sample_count_r\[6\] _1007_ VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_4_52 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3113_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0013_ net93 core.cnb.shift_register_r\[11\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA__2448__B1 core.pdc.rowon_bottotop_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3044_ VSS VDD _0930_ _0932_ _0918_ VSS VDD sky130_fd_sc_hd__nand2_1
Xgenblk1\[4\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[4\] core.pdc.col_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2828_ VSS VDD _0723_ _0644_ _0679_ _0722_ VSS VDD sky130_fd_sc_hd__and3_1
X_2759_ VSS VDD _0649_ _0652_ _0655_ _0654_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_86_464 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_328 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_339 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_86_486 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_fanout57_A net58 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1662__A1 _1199_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout73 VSS VDD net83 net73 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout62 VDD VSS net62 net63 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout84 VSS VDD net85 net84 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_80_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_61 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[6\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[6\] core.ndc.row_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_49_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_412 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_309 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_489 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1992_ VSS VDD _1082_ _1114_ _0087_ _1412_ VSS VDD sky130_fd_sc_hd__o21ai_2
X_2613_ VSS VDD _0519_ core.osr.next_result_w\[2\] core.osr.next_result_w\[4\] _1003_
+ _0523_ _0520_ VSS VDD sky130_fd_sc_hd__o221a_1
XFILLER_133_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2544_ VDD VSS _0466_ _0465_ _0467_ _0468_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_2475_ VSS VDD core.pdc.row_out_n\[7\] core.pdc.rowoff_out_n\[7\] core.pdc.rowon_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1426_ VDD VSS _0990_ core.osr.osr_mode_r\[1\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_83_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_467 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3027_ VDD VSS _0915_ _0914_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_83_489 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_132_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[1\].buf_n_coln VDD VSS core.ndc.col_out_n\[1\] nmatrix_col_core_n_buffered\[1\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_115_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3181__RESET_B net86 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2260_ VDD VSS core.osr.next_result_w\[5\] _0288_ VSS VDD sky130_fd_sc_hd__inv_2
X_2191_ VDD VSS _0228_ _0227_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_37_136 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[0] nmatrix_col_core_n_buffered\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_92_275 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_92_286 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1975_ VSS VDD _0074_ _1141_ _1389_ _1111_ VSS VDD sky130_fd_sc_hd__mux2_1
Xpmat pmatrix_row_core_n_buffered\[0\] pmatrix_row_core_n_buffered\[1\] pmatrix_row_core_n_buffered\[2\]
+ pmatrix_row_core_n_buffered\[3\] pmatrix_row_core_n_buffered\[4\] pmatrix_row_core_n_buffered\[5\]
+ pmatrix_row_core_n_buffered\[6\] pmatrix_row_core_n_buffered\[7\] pmatrix_row_core_n_buffered\[8\]
+ pmatrix_row_core_n_buffered\[9\] pmatrix_row_core_n_buffered\[10\] pmatrix_row_core_n_buffered\[11\]
+ pmatrix_row_core_n_buffered\[12\] pmatrix_row_core_n_buffered\[13\] pmatrix_row_core_n_buffered\[14\]
+ pmatrix_row_core_n_buffered\[15\] pmatrix_rowon_core_n_buffered\[0\] pmatrix_rowon_core_n_buffered\[1\]
+ pmatrix_rowon_core_n_buffered\[2\] pmatrix_rowon_core_n_buffered\[3\] pmatrix_rowon_core_n_buffered\[4\]
+ pmatrix_rowon_core_n_buffered\[5\] pmatrix_rowon_core_n_buffered\[6\] pmatrix_rowon_core_n_buffered\[7\]
+ pmatrix_rowon_core_n_buffered\[8\] pmatrix_rowon_core_n_buffered\[9\] pmatrix_rowon_core_n_buffered\[10\]
+ pmatrix_rowon_core_n_buffered\[11\] pmatrix_rowon_core_n_buffered\[12\] pmatrix_rowon_core_n_buffered\[13\]
+ pmatrix_rowon_core_n_buffered\[14\] pmatrix_rowon_core_n_buffered\[15\] core.pdc.rowoff_out_n\[0\]
+ core.pdc.rowoff_out_n\[1\] core.pdc.rowoff_out_n\[2\] core.pdc.rowoff_out_n\[3\]
+ core.pdc.rowoff_out_n\[4\] core.pdc.rowoff_out_n\[5\] core.pdc.rowoff_out_n\[6\]
+ core.pdc.rowoff_out_n\[7\] core.pdc.rowoff_out_n\[8\] core.pdc.rowoff_out_n\[9\]
+ core.pdc.rowoff_out_n\[10\] core.pdc.rowoff_out_n\[11\] core.pdc.rowoff_out_n\[12\]
+ core.pdc.rowoff_out_n\[13\] core.pdc.rowoff_out_n\[14\] core.pdc.rowoff_out_n\[15\]
+ vcm/vcm sample_pmatrix_cgen _0000_ pmatrix_col_core_n_buffered\[31\] pmatrix_col_core_n_buffered\[30\]
+ pmatrix_col_core_n_buffered\[29\] pmatrix_col_core_n_buffered\[28\] pmatrix_col_core_n_buffered\[27\]
+ pmatrix_col_core_n_buffered\[26\] pmatrix_col_core_n_buffered\[25\] pmatrix_col_core_n_buffered\[24\]
+ pmatrix_col_core_n_buffered\[23\] pmatrix_col_core_n_buffered\[22\] pmatrix_col_core_n_buffered\[21\]
+ pmatrix_col_core_n_buffered\[20\] pmatrix_col_core_n_buffered\[19\] pmatrix_col_core_n_buffered\[18\]
+ pmatrix_col_core_n_buffered\[17\] pmatrix_col_core_n_buffered\[16\] pmatrix_col_core_n_buffered\[15\]
+ pmatrix_col_core_n_buffered\[14\] pmatrix_col_core_n_buffered\[13\] pmatrix_col_core_n_buffered\[12\]
+ pmatrix_col_core_n_buffered\[11\] pmatrix_col_core_n_buffered\[10\] pmatrix_col_core_n_buffered\[9\]
+ pmatrix_col_core_n_buffered\[8\] pmatrix_col_core_n_buffered\[7\] pmatrix_col_core_n_buffered\[6\]
+ pmatrix_col_core_n_buffered\[5\] pmatrix_col_core_n_buffered\[4\] pmatrix_col_core_n_buffered\[3\]
+ pmatrix_col_core_n_buffered\[2\] pmatrix_col_core_n_buffered\[1\] pmatrix_col_core_n_buffered\[0\]
+ core.cnb.data_register_r\[2\] core.cnb.data_register_r\[1\] core.cnb.data_register_r\[0\]
+ net95 pmat_sample_switch_buffered pmat_sample_switch_n_buffered inp_analog core.pdc.col_out\[0\]
+ core.pdc.col_out\[1\] core.pdc.col_out\[2\] core.pdc.col_out\[3\] core.pdc.col_out\[4\]
+ core.pdc.col_out\[5\] core.pdc.col_out\[6\] core.pdc.col_out\[7\] core.pdc.col_out\[8\]
+ core.pdc.col_out\[9\] core.pdc.col_out\[10\] core.pdc.col_out\[11\] core.pdc.col_out\[12\]
+ core.pdc.col_out\[13\] core.pdc.col_out\[14\] core.pdc.col_out\[15\] core.pdc.col_out\[16\]
+ core.pdc.col_out\[17\] core.pdc.col_out\[18\] core.pdc.col_out\[19\] core.pdc.col_out\[20\]
+ core.pdc.col_out\[21\] core.pdc.col_out\[22\] core.pdc.col_out\[23\] core.pdc.col_out\[24\]
+ core.pdc.col_out\[25\] core.pdc.col_out\[26\] core.pdc.col_out\[27\] core.pdc.col_out\[28\]
+ core.pdc.col_out\[29\] core.pdc.col_out\[30\] core.pdc.col_out\[31\] ctop_pmatrix_analog
+ VSS VDD adc_array_matrix_12bit
XFILLER_20_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_106_119 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3174__CLK net58 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col[16] core.ndc.col_out\[16\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2527_ VSS VDD _0017_ _0455_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_88_515 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2458_ VSS VDD core.ndc.row_out_n\[3\] core.ndc.rowoff_out_n\[3\] core.ndc.rowon_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2389_ VSS VDD _0985_ _0397_ _0401_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_28_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_56_489 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1502__A _1053_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2317__B core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_62 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_120_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_136 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2243__A core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1760_ VSS VDD _1274_ _1131_ _1243_ VSS VDD sky130_fd_sc_hd__or2_1
X_1691_ VSS VDD _1035_ _1225_ _1153_ _1224_ core.ndc.col_out_n\[12\] _1226_ VSS VDD
+ sky130_fd_sc_hd__o221a_2
X_2312_ VSS VDD _0251_ _0336_ _0335_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_111_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2243_ VSS VDD core.cnb.result_out\[4\] _0273_ core.osr.result_r\[4\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2174_ VDD VSS _0214_ _0193_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_cgen_dlycontrol4_in[4] net7 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1958_ VSS VDD _1047_ _1057_ _1410_ _1409_ VSS VDD sky130_fd_sc_hd__o21ai_2
X_1889_ VSS VDD _1306_ _1362_ core.pdc.rowon_out_n\[1\] _1364_ VSS VDD sky130_fd_sc_hd__o21ai_2
Xoutput39 VDD VSS result_out[10] net39 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_102_111 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1550__A3 _1105_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_56_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_128 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_42 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2047__B _1235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_col[2] core.pdc.col_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_43 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[9\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[9\] core.pdc.col_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_90_510 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2930_ VSS VDD _0638_ _0766_ _0822_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_15_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2861_ VSS VDD _0691_ _0756_ _0208_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1812_ VDD VSS _1305_ _1304_ VSS VDD sky130_fd_sc_hd__inv_2
X_2792_ VSS VDD _0208_ _0688_ _0670_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1743_ VSS VDD _1265_ _1227_ _1225_ VSS VDD sky130_fd_sc_hd__or2_1
X_1674_ VSS VDD _1212_ _1214_ _1213_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_97_131 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2226_ VDD VSS _0258_ _0256_ _0257_ VSS VDD sky130_fd_sc_hd__and2_1
X_2157_ VSS VDD _0201_ core.cnb.average_counter_r\[4\] _0187_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_26_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2493__A1 core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2088_ VSS VDD _1227_ _0072_ _0151_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_13_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_fanout87_A net94 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_67_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_123_96 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_83_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_genblk1\[14\].buf_n_coln_A core.ndc.col_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[17] nmatrix_col_core_n_buffered\[17\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3060_ VSS VDD _0945_ _0947_ _0507_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2011_ VSS VDD _0101_ _0102_ _1275_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_90_340 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_237 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2913_ VDD VSS _0805_ _0804_ VSS VDD sky130_fd_sc_hd__inv_2
X_2844_ VDD VSS _0739_ core.cnb.shift_register_r\[11\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1738__B1 _1035_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2775_ VSS VDD core.cnb.shift_register_r\[16\] _0670_ _0671_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1726_ VSS VDD _1254_ _1253_ _1252_ _1250_ VSS VDD sky130_fd_sc_hd__and3_1
X_1657_ VDD VSS _1052_ _1199_ _1059_ _1036_ VSS VDD sky130_fd_sc_hd__o21ai_4
X_1588_ VSS VDD _1138_ _1137_ _1077_ _1133_ VSS VDD sky130_fd_sc_hd__mux2_1
Xgenblk1\[6\].buf_n_coln VDD VSS core.ndc.col_out_n\[6\] nmatrix_col_core_n_buffered\[6\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_2209_ VDD VSS _0239_ core.osr.next_result_w\[0\] _0242_ VSS VDD sky130_fd_sc_hd__xor2_1
X_3189_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0059_ net81 core.cnb.data_register_r\[9\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA__3108__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1510__A _1047_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2325__B _0255_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_118_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_118_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_78_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_440 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_89_473 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_94_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1968__B1 _1088_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2251__A core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2560_ VSS VDD core.cnb.data_register_r\[2\] _0482_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2491_ VDD VSS net17 _1040_ net16 _0436_ VSS VDD sky130_fd_sc_hd__or3_1
X_1511_ VSS VDD _1068_ _1069_ _1037_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1442_ VSS VDD _1006_ _1005_ _0998_ _0997_ _0988_ VSS VDD sky130_fd_sc_hd__and4_1
XFILLER_4_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__3082__A _0758_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3112_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0012_ net93 core.cnb.shift_register_r\[10\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3043_ VDD VSS _0831_ _0930_ _0856_ _0931_ VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_139_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2827_ VDD VSS _0722_ _0659_ VSS VDD sky130_fd_sc_hd__inv_2
X_2758_ VSS VDD core.cnb.shift_register_r\[11\] _0653_ _0654_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1709_ VSS VDD _1240_ _1241_ _1213_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2689_ VSS VDD core.osr.next_result_w\[13\] _0590_ _0535_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1505__A core.ndc.col_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_498 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout74 VDD VSS net74 net76 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout63 VDD VSS net63 net66 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout85 VDD VSS net85 net87 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_13_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_89_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2071__A _0081_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_178 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1991_ VDD VSS core.pdc.col_out_n\[6\] core.pdc.col_out\[6\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__2602__A1 core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2612_ VDD VSS _0521_ net45 _0395_ _0035_ _0522_ VSS VDD sky130_fd_sc_hd__a22o_1
X_2543_ VSS VDD _0181_ _0207_ _0467_ core.cnb.average_sum_r\[1\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_2474_ VSS VDD core.pdc.rowon_out_n\[6\] core.pdc.rowoff_out_n\[6\] core.pdc.row_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1425_ VDD VSS _0989_ core.osr.osr_mode_r\[0\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_18_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1979__B _1155_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3026_ VSS VDD _0475_ _0914_ _0913_ _1117_ _0911_ VSS VDD sky130_fd_sc_hd__o211ai_1
XFILLER_34_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_310 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_91_490 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_398 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xnmat_sample_buf_n VSS VDD nmat_sample_switch_n_buffered core.cnb.enable_loop_out
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1995__A _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_59_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_132_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_132_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_75_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_75_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_131_30 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2190_ VSS VDD _0226_ _0223_ _0227_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_1_21 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1974_ VDD VSS core.pdc.col_out\[4\] core.pdc.col_out_n\[4\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_136_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_114_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col[15] core.ndc.col_out\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2526_ VSS VDD _0455_ _0454_ _0219_ core.cnb.shift_register_r\[15\] VSS VDD sky130_fd_sc_hd__mux2_1
X_2457_ VSS VDD core.ndc.row_out_n\[2\] core.ndc.rowoff_out_n\[2\] core.ndc.rowon_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_29_17 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2388_ VSS VDD core.osr.sample_count_r\[2\] _0398_ _0400_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_45_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3009_ VSS VDD _0884_ _0877_ _0898_ _0895_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_10_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_126_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_126_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_120_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__3058__A1 _0799_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_35_82 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1690_ VSS VDD _1172_ _1226_ _1093_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1792__B2 _1125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2897__C _1395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2311_ VDD VSS _0335_ core.cnb.result_out\[10\] VSS VDD sky130_fd_sc_hd__inv_2
X_2242_ VSS VDD _0272_ core.cnb.result_out\[4\] core.osr.result_r\[4\] VSS VDD sky130_fd_sc_hd__or2_1
X_2173_ VSS VDD core.cnb.next_average_counter_w\[3\] _0213_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1603__A core.ndc.col_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2137__C core.cnb.sampled_avg_control_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol4_in[3] net6 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3141__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1957_ VDD VSS _1409_ _1400_ VSS VDD sky130_fd_sc_hd__buf_2
X_1888_ VSS VDD _1363_ _1364_ _1303_ VSS VDD sky130_fd_sc_hd__nor2_2
X_2509_ VSS VDD _0446_ core.cnb.shift_register_r\[8\] _0444_ core.cnb.shift_register_r\[7\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_102_123 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1513__A core.cnb.data_register_r\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[2\].buf_p_rown_A core.pdc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_54 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_98 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_522 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2860_ VSS VDD _0718_ _0754_ _0755_ _0719_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1811_ VSS VDD _1303_ _1304_ core.cnb.data_register_r\[10\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2791_ VSS VDD _0686_ _0687_ core.cnb.data_register_r\[0\] VSS VDD sky130_fd_sc_hd__nand2_1
X_1742_ VDD VSS _1263_ _1264_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_1673_ VDD VSS _1213_ _1092_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_97_143 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2225_ VSS VDD core.cnb.result_out\[2\] _0257_ core.osr.result_r\[2\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2429__A _1342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2156_ VSS VDD _0193_ _0196_ _0200_ _0199_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_26_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2493__A2 _0220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_235 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_246 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_393 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2087_ VDD VSS core.pdc.col_out\[22\] core.pdc.col_out_n\[22\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA_nmat_sample_buf_A net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2989_ VSS VDD _0877_ _0879_ _0878_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_123_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__3187__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[12\].buf_p_rowonn_A core.pdc.rowon_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[4] net23 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[16] nmatrix_col_core_n_buffered\[16\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2010_ VSS VDD _0101_ _1085_ _1395_ _1390_ _1132_ VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_76_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1600__B _1032_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2912_ VSS VDD _0802_ _0804_ _0803_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2843_ VSS VDD _0732_ _0734_ _0738_ _0737_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2774_ VSS VDD _0637_ _0670_ VSS VDD sky130_fd_sc_hd__inv_1
XANTENNA__1738__A1 _1259_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1725_ VSS VDD _1182_ _1253_ _1177_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1656_ VSS VDD _1198_ _1186_ _1054_ _1197_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1587_ VSS VDD _1122_ _1137_ _1136_ VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_85_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2208_ VSS VDD _0241_ _0242_ core.osr.result_r\[0\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_67_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3188_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0058_ net87 core.cnb.data_register_r\[8\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_4
X_2139_ VSS VDD _0181_ _0183_ _0182_ VSS VDD sky130_fd_sc_hd__nand2_1
Xgenblk2\[3\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[3\] core.pdc.rowon_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_139_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_118_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_118_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_134_52 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_89_485 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_134_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_94_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_input12_A config_1_in[4] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1701__A net15 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_43_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2490_ VDD VSS net36 _0435_ VSS VDD sky130_fd_sc_hd__inv_2
X_1510_ VDD VSS _1068_ _1047_ VSS VDD sky130_fd_sc_hd__inv_2
X_1441_ VSS VDD core.osr.sample_count_r\[6\] _1003_ _1001_ _0999_ _1005_ _1004_ VSS
+ VDD sky130_fd_sc_hd__o221a_1
X_3111_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0011_ net90 core.cnb.shift_register_r\[9\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_67_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_3042_ VSS VDD _0930_ _0910_ _0833_ _0726_ _0929_ VSS VDD sky130_fd_sc_hd__and4_1
XANTENNA__1656__A0 _1197_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_382 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_182 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_23_19 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_sample_buf_n_A core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2442__A core.ndc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2826_ VDD VSS _0719_ _0718_ _0720_ _0721_ VSS VDD sky130_fd_sc_hd__a21o_1
X_2757_ VDD VSS _0653_ core.cnb.shift_register_r\[10\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_2_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2688_ VSS VDD _0347_ _0568_ _0589_ _0348_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1708_ VDD VSS _1240_ _1108_ VSS VDD sky130_fd_sc_hd__inv_2
X_1639_ VDD VSS _1183_ _1182_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_input4_A config_1_in[11] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_411 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_86_444 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_104_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xfanout64 VSS VDD net66 net64 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout75 VDD VSS net75 net76 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout86 VDD VSS net86 net87 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2071__B _1213_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_clk_dig_dummy_A clknet_0_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_127 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1990_ VSS VDD _0086_ core.pdc.col_out_n\[6\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__2262__A core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_118_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2611_ VSS VDD _0288_ _0522_ _0517_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2542_ VDD VSS core.cnb.average_sum_r\[2\] _0195_ _0198_ _0466_ VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA_nmat_col[31] core.ndc.col_out\[31\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3093__A _0758_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2473_ VSS VDD core.pdc.row_out_n\[4\] core.pdc.rowoff_out_n\[4\] core.pdc.rowon_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1424_ VSS VDD _0987_ _0988_ _0983_ VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_83_414 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1629__B1 _1118_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_127 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3025_ VSS VDD _0912_ _0472_ _0913_ _0911_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__2172__A _0210_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2809_ VDD VSS _0704_ _0703_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_117_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_115_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_131_42 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_61_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_91_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xnmat_96 nmat_96/LO net96 VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__3190__RESET_B net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xcomp comp/clk ctop_pmatrix_analog ctop_nmatrix_analog decision_finish_comp_n comp/latch_qn
+ core.cnb.comparator_in VDD VSS VSS adc_comp_latch
XFILLER_37_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_92_200 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1973_ VDD VSS _1121_ _0068_ core.pdc.col_out\[4\] _0070_ _1296_ _0073_ VSS VDD sky130_fd_sc_hd__a221o_1
XFILLER_60_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col[14] core.ndc.col_out\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2525_ VSS VDD core.cnb.shift_register_r\[16\] _0454_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2456_ VSS VDD core.ndc.rowon_out_n\[1\] core.ndc.rowoff_out_n\[1\] core.ndc.row_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_29_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2387_ VDD VSS core.osr.next_sample_count_w\[1\] _0399_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_83_211 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2167__A _0210_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3008_ VSS VDD _0887_ _0897_ _0896_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_299 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_73 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3191__SET_B net82 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_469 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_491 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_42_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1792__A2 _1279_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2310_ VSS VDD _0331_ _0255_ _0334_ _0333_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2241_ VSS VDD _0988_ _0271_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_111_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2172_ VSS VDD _0213_ _0193_ _0194_ _0210_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_46_491 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_cgen_dlycontrol4_in[2] net5 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1956_ VDD VSS core.pdc.col_out_n\[2\] core.pdc.col_out\[2\] VSS VDD sky130_fd_sc_hd__inv_2
X_1887_ VDD VSS _1363_ _1029_ VSS VDD sky130_fd_sc_hd__inv_2
X_2508_ VSS VDD _0008_ _0445_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_102_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1940__C1 _1085_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2439_ VSS VDD _1376_ core.ndc.rowon_out_n\[2\] _1385_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_56_255 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_112_66 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_24_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_21_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_62_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1810_ VSS VDD core.cnb.data_register_r\[9\] _1303_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_7_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2790_ VSS VDD _0677_ _0685_ _0686_ VSS VDD sky130_fd_sc_hd__nand2b_1
X_1741_ VSS VDD _1033_ _1153_ _1263_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2270__A core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1672_ VDD VSS _1207_ _1103_ _1206_ _1212_ VSS VDD sky130_fd_sc_hd__a21o_1
X_2224_ VSS VDD _0256_ core.cnb.result_out\[2\] core.osr.result_r\[2\] VSS VDD sky130_fd_sc_hd__or2_1
X_2155_ VSS VDD _0197_ _0198_ _0199_ core.cnb.average_counter_r\[3\] VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_93_361 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2086_ VDD VSS _0101_ _1173_ core.pdc.col_out\[22\] _0103_ _1096_ _0150_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2988_ VSS VDD _0874_ _1113_ _0878_ _0875_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1939_ VDD VSS core.cnb.data_register_r\[3\] _1395_ VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__2180__A _0208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_16_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[15\].buf_p_rown_A core.pdc.row_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[3] net22 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3131__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[15] nmatrix_col_core_n_buffered\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2911_ VSS VDD _0798_ _1200_ _0803_ _0800_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2842_ VSS VDD _0736_ _0725_ _0737_ _0724_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2773_ VSS VDD _0669_ _0635_ _0206_ _0668_ VSS VDD sky130_fd_sc_hd__and3_1
X_1724_ VSS VDD _1251_ _1252_ _1213_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1655_ VDD VSS _1196_ _1197_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_1586_ VDD VSS _1136_ _1135_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_85_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2207_ VSS VDD _0240_ _0241_ VSS VDD sky130_fd_sc_hd__clkbuf_4
X_3187_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0057_ net85 core.cnb.data_register_r\[7\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_4
X_2138_ VSS VDD _0182_ core.cnb.average_counter_r\[1\] core.cnb.average_counter_r\[0\]
+ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1998__B _1155_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2069_ VSS VDD _1075_ _0115_ _0069_ _1126_ core.pdc.col_out_n\[18\] _0141_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout92_A net94 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_497 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_94_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_134_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_94_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_94_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_84 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1968__A2 _1104_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1440_ VSS VDD _1004_ core.osr.sample_count_r\[8\] _0992_ VSS VDD sky130_fd_sc_hd__or2_1
X_3110_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0010_ net90 core.cnb.shift_register_r\[8\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA_genblk1\[10\].buf_n_coln_A core.ndc.col_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3041_ VSS VDD _0929_ _0818_ _0827_ _0745_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__1656__A1 _1186_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2605__B1 _0395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2825_ VDD VSS _0720_ _0687_ VSS VDD sky130_fd_sc_hd__inv_2
X_2756_ VSS VDD _0651_ _0646_ _0652_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2687_ VDD VSS _1008_ _0376_ _0524_ _0588_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_1707_ VDD VSS _1238_ _1239_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_1638_ VSS VDD _1061_ _1182_ _1053_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1569_ VDD VSS _1121_ _1101_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_46_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_104_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_104_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_104_45 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[12\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[12\] core.pdc.row_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2617__B _1002_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_120_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xfanout65 VSS VDD net65 net66 VSS VDD sky130_fd_sc_hd__clkbuf_1
Xfanout54 VDD VSS net54 net55 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA_cgen_dlycontrol2_in[4] net33 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_42 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout76 VSS VDD net82 net76 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout87 VDD VSS net87 net94 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_80_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_86 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_89_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_158 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_92_404 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1712__A _1034_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2610_ VSS VDD _0521_ _0517_ core.osr.next_result_w\[3\] _0519_ _0520_ VSS VDD sky130_fd_sc_hd__o211a_1
X_2541_ VSS VDD _0462_ _0463_ _0465_ _0464_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_126_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2472_ VSS VDD core.pdc.row_out_n\[3\] core.pdc.rowoff_out_n\[3\] core.pdc.rowon_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1423_ VSS VDD _0987_ _0986_ _0985_ core.osr.sample_count_r\[0\] _0984_ VSS VDD sky130_fd_sc_hd__and4b_1
XANTENNA__1629__A1 _1085_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_139 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3024_ VSS VDD _0835_ _0834_ _0912_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2437__B core.pdc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2808_ VSS VDD _0674_ _0703_ _0702_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2739_ VSS VDD core.cnb.shift_register_r\[6\] core.cnb.shift_register_r\[7\] _0635_
+ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1565__A0 _1112_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_86_253 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2347__B _0240_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_108_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1588__S _1077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1972_ VSS VDD _0065_ _0072_ _0073_ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk2\[12\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[12\] core.ndc.rowon_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA_nmat_col[13] core.ndc.col_out\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2524_ VSS VDD _0016_ _0453_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2455_ VSS VDD core.pdc.rowon_out_n\[0\] _1362_ core.ndc.rowon_out_n\[14\] _1365_
+ VSS VDD sky130_fd_sc_hd__o21ai_2
X_2386_ VDD VSS _0398_ core.osr.is_last_sample _0396_ _0399_ VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_28_106 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_45_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3007_ VSS VDD _0895_ _0896_ VSS VDD sky130_fd_sc_hd__clkinvlp_2
XANTENNA__2183__A core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_101_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_124_7 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_144 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_42_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2240_ VSS VDD _0270_ core.osr.next_result_w\[3\] VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2171_ VSS VDD core.cnb.next_average_counter_w\[2\] _0212_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA_cgen_dlycontrol4_in[1] net4 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[13\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[13\] core.pdc.col_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1955_ VDD VSS _1398_ _1279_ core.pdc.col_out\[2\] _1406_ _1296_ _1408_ VSS VDD sky130_fd_sc_hd__a221o_1
X_1886_ VSS VDD _1038_ _1362_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2507_ VSS VDD _0445_ core.cnb.shift_register_r\[7\] _0444_ core.cnb.shift_register_r\[6\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__1940__B1 _1079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2438_ VDD VSS _1340_ _1027_ _1364_ core.ndc.rowon_out_n\[1\] VSS VDD sky130_fd_sc_hd__a21o_1
X_2369_ VDD VSS _0386_ _0381_ _0385_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_112_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_112_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_115_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_97_24 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col_n[31] nmatrix_col_core_n_buffered\[31\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input35_A start_conversion_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2088__A _1227_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1720__A core.ndc.col_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_62_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1740_ VSS VDD _1157_ _1262_ _1152_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_7_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1671_ VDD VSS _1210_ _1211_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_2223_ VSS VDD _0988_ _0255_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2154_ VDD VSS _0198_ _0181_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_16_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1630__A _1175_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2085_ VDD VSS _0150_ _0149_ VSS VDD sky130_fd_sc_hd__inv_2
Xgenblk2\[9\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[9\] core.ndc.rowon_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2987_ VSS VDD _0876_ _0877_ _1058_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2461__A core.ndc.row_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1938_ VDD VSS _1394_ _1388_ VSS VDD sky130_fd_sc_hd__buf_2
X_1869_ VSS VDD net14 _1308_ _1351_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_123_11 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_123_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk1\[10\].buf_n_coln VDD VSS core.ndc.col_out_n\[10\] nmatrix_col_core_n_buffered\[10\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__1540__A _1095_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_16_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_281 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_32_52 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2090__B _1235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1715__A core.ndc.col_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[2] net21 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[14] nmatrix_col_core_n_buffered\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2910_ VSS VDD _0801_ _0802_ _1055_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2841_ VSS VDD _0646_ _0735_ _0736_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2772_ VSS VDD core.cnb.shift_register_r\[2\] _0667_ _0668_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1723_ VDD VSS _1251_ _1049_ VSS VDD sky130_fd_sc_hd__inv_2
X_1654_ VSS VDD _1195_ _1196_ _1051_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1585_ VSS VDD _1135_ _1134_ _1050_ VSS VDD sky130_fd_sc_hd__nor2_4
X_2206_ VDD VSS _0240_ _0988_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_54_502 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3186_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0056_ net85 core.cnb.data_register_r\[6\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_2137_ VSS VDD _0176_ _0180_ _0181_ core.cnb.sampled_avg_control_r\[0\] VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__2456__A core.ndc.rowon_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2068_ VSS VDD _0120_ _0141_ _1155_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_5_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_118_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1535__A _1092_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_134_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout85_A net87 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_94_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk2\[14\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[14\] core.ndc.row_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_27_63 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1968__A3 _1105_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3184__RESET_B net87 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_67 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3040_ VSS VDD _0926_ _1055_ _0928_ _0927_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_51_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2824_ VSS VDD _0714_ _0716_ _0719_ core.cnb.pswitch_out\[1\] VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_136_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2755_ VSS VDD _0650_ _0651_ _0642_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2686_ VSS VDD _0585_ _0044_ _0587_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1706_ VSS VDD _1227_ _1166_ _1238_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1637_ VSS VDD _1180_ _1181_ _1096_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1568_ VDD VSS core.ndc.col_out\[3\] core.ndc.col_out_n\[3\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_48_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_86_424 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_58_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1499_ VSS VDD _1059_ _1058_ _1044_ VSS VDD sky130_fd_sc_hd__nand2_2
X_3169_ VSS VDD net66 core.osr.next_result_w\[9\] net76 core.osr.result_r\[9\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_104_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_398 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_120_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2633__B core.osr.next_result_w\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout55 VSS VDD core.cnb.is_sampling_w net55 VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_80_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_cgen_dlycontrol2_in[3] net32 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout88 VSS VDD net92 net88 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout77 VDD VSS net77 net80 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout66 VSS VDD net67 net66 VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__3121__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_129_76 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_98 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2532__A0 core.cnb.sampled_avg_control_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_295 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_38_62 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1712__B _1243_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[18\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[18\] core.pdc.col_out_n\[18\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_118_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2540_ VSS VDD _0231_ _0177_ _0464_ _0186_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_2471_ VSS VDD core.pdc.row_out_n\[2\] core.pdc.rowoff_out_n\[2\] core.pdc.rowon_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1422_ VSS VDD core.osr.sample_count_r\[5\] core.osr.sample_count_r\[3\] core.osr.sample_count_r\[1\]
+ _0986_ VSS VDD sky130_fd_sc_hd__nor3_1
XANTENNA__1903__A _1342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3023_ VSS VDD _0910_ _0911_ _0827_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_346 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2807_ VSS VDD _0702_ _0639_ _0701_ _0699_ VSS VDD sky130_fd_sc_hd__nand3b_1
X_2738_ VSS VDD _0633_ _0634_ core.cnb.shift_register_r\[9\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1565__A1 _1118_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2669_ VDD VSS _0565_ _0572_ _0042_ _0571_ VSS VDD sky130_fd_sc_hd__o21bai_1
Xgenblk1\[20\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[20\] core.pdc.col_out_n\[20\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_86_265 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2644__A core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_37 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_64 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_40_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_108_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3167__CLK net61 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_65_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2554__A core.cnb.pswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1971_ VDD VSS _0072_ _0071_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col[12] core.ndc.col_out\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2523_ VSS VDD _0453_ core.cnb.shift_register_r\[15\] _0219_ core.cnb.shift_register_r\[14\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_46_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2454_ VDD VSS core.ndc.rowon_out_n\[13\] _0431_ VSS VDD sky130_fd_sc_hd__inv_2
X_2385_ VDD VSS _0398_ _0397_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_cgen_dlycontrol1_in[4] net28 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_28_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput1 VSS VDD net1 clk_vcm VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_56_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[15\].buf_n_coln VDD VSS core.ndc.col_out_n\[15\] nmatrix_col_core_n_buffered\[15\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_3006_ VSS VDD _0893_ _0895_ _0894_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_10_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_111_126 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2170_ VSS VDD _0212_ _0197_ _0192_ _0210_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__1900__B _1022_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol4_in[0] net3 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1954_ VSS VDD _1272_ _1407_ _1408_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1885_ VSS VDD core.pdc.row_out_n\[15\] _1361_ core.ndc.rowon_out_n\[0\] VSS VDD
+ sky130_fd_sc_hd__nand2_2
X_2506_ VSS VDD _0208_ _0444_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_88_316 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2437_ VSS VDD _1341_ core.ndc.row_out_n\[15\] core.pdc.rowon_out_n\[0\] VSS VDD
+ sky130_fd_sc_hd__nand2_1
X_2368_ VDD VSS _0385_ _0384_ _0255_ VSS VDD sky130_fd_sc_hd__and2_1
X_2299_ VSS VDD _0309_ _0307_ _0323_ _0317_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_24_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1538__A core.ndc.col_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2641__B core.osr.next_result_w\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2088__B _0072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3138__RESET_B net85 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input28_A config_2_in[4] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_34 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1670_ VSS VDD _1033_ _1209_ _1210_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2222_ VDD VSS core.osr.next_result_w\[1\] _0254_ VSS VDD sky130_fd_sc_hd__inv_2
X_2153_ VSS VDD _0191_ _0197_ _0184_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_53_216 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2084_ VSS VDD _0149_ _1039_ _0113_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_21_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_21_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_124 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2986_ VSS VDD _0874_ _0876_ _0875_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1937_ VDD VSS core.pdc.col_out_n\[0\] core.pdc.col_out\[0\] VSS VDD sky130_fd_sc_hd__inv_2
X_1868_ VSS VDD _1324_ _1333_ _1350_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1799_ VDD VSS _1121_ _1083_ core.ndc.col_out\[30\] _1247_ _1296_ _1298_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_88_168 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_123_23 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_396 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_293 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_146 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_cgen_dlycontrol3_in[1] net20 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[13] nmatrix_col_core_n_buffered\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_87_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_300 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_208 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2840_ VSS VDD _0663_ _0735_ _0641_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2771_ VDD VSS _0667_ core.cnb.shift_register_r\[3\] VSS VDD sky130_fd_sc_hd__inv_2
X_1722_ VSS VDD _1249_ _1250_ _1102_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1653_ VSS VDD _1066_ _1195_ _1104_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1584_ VSS VDD core.cnb.data_register_r\[6\] core.cnb.data_register_r\[5\] _1134_
+ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk1\[25\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[25\] core.pdc.col_out_n\[25\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2205_ VDD VSS _0239_ core.cnb.result_out\[0\] VSS VDD sky130_fd_sc_hd__inv_2
X_3185_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0055_ net87 core.cnb.data_register_r\[5\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2136_ VDD VSS _0180_ core.cnb.sampled_avg_control_r\[2\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2456__B core.ndc.row_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_514 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2067_ VDD VSS core.pdc.col_out\[17\] core.pdc.col_out_n\[17\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2969_ VSS VDD _0861_ _0805_ _0860_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1551__A _1106_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_182 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2382__A _0395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_rowoff_n[8] core.pdc.rowoff_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1461__A _1022_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2557__A _0438_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_374 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_90_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2066__B1 _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2605__A2 _0995_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2823_ VSS VDD _0717_ _0718_ core.cnb.data_register_r\[1\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_76_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2754_ VSS VDD core.cnb.shift_register_r\[8\] core.cnb.shift_register_r\[9\] _0650_
+ VSS VDD sky130_fd_sc_hd__nor2_1
X_1705_ VDD VSS core.ndc.col_out\[13\] core.ndc.col_out_n\[13\] VSS VDD sky130_fd_sc_hd__inv_2
X_2685_ VDD VSS _0587_ _0586_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1636__A _1129_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1636_ VDD VSS _1180_ _1129_ VSS VDD sky130_fd_sc_hd__inv_2
X_1567_ VSS VDD _1075_ _1109_ _1108_ _1064_ core.ndc.col_out_n\[3\] _1120_ VSS VDD
+ sky130_fd_sc_hd__o221a_2
X_1498_ VSS VDD core.cnb.data_register_r\[6\] _1058_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_86_436 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3168_ VSS VDD net66 core.osr.next_result_w\[8\] net76 core.osr.result_r\[8\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_104_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2119_ VSS VDD core.pdc.col_out_n\[29\] _0169_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_3099_ VSS VDD _0981_ core.osr.osr_mode_r\[2\] _0241_ net13 VSS VDD sky130_fd_sc_hd__mux2_1
Xfanout56 VDD VSS net56 net57 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cgen_dlycontrol2_in[2] net31 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout89 VDD VSS net89 net92 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout78 VDD VSS net78 net80 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout67 VSS VDD net37 net67 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_129_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1546__A _1101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[22\].buf_n_coln VDD VSS core.ndc.col_out_n\[22\] nmatrix_col_core_n_buffered\[22\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_49_116 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_38_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_428 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input10_A config_1_in[2] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_61 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1456__A _0983_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2470_ VSS VDD core.pdc.row_out_n\[1\] core.pdc.rowoff_out_n\[1\] core.pdc.rowon_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1421_ VDD VSS _0985_ core.osr.sample_count_r\[2\] VSS VDD sky130_fd_sc_hd__inv_2
X_3022_ VDD VSS _0910_ _0809_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_63_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2806_ VSS VDD _0700_ _0659_ _0701_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2737_ VDD VSS _0633_ core.cnb.shift_register_r\[8\] VSS VDD sky130_fd_sc_hd__inv_2
X_2668_ VDD VSS _0394_ core.osr.next_result_w\[4\] _0542_ _0572_ net52 VSS VDD sky130_fd_sc_hd__a22o_1
X_1619_ VSS VDD _1165_ _1164_ _1041_ _1161_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_59_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2599_ VDD VSS _0439_ _0335_ _0512_ _0032_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_115_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input2_A config_1_in[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_17 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2644__B _1002_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_24_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_138_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_40_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_123_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1970_ VSS VDD _0071_ _1115_ _1052_ _1389_ _1045_ VSS VDD sky130_fd_sc_hd__a31o_1
X_2522_ VSS VDD _0015_ _0452_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2453_ VSS VDD _1380_ _0431_ _1306_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_sample_p_in net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2384_ VSS VDD core.osr.sample_count_r\[0\] _0397_ core.osr.sample_count_r\[1\] VSS
+ VDD sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_dlycontrol1_in[3] net27 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput2 VSS VDD net2 config_1_in[0] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__3111__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3005_ VSS VDD _0890_ _1051_ _0894_ _0891_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_36_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2480__A core.pdc.rowon_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_105_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_21 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout60_A net61 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_439 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1718__B _1093_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1734__A core.ndc.col_out_n\[17\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3134__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2549__B _0438_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1953_ VSS VDD _1123_ _1403_ _1068_ _1407_ VSS VDD sky130_fd_sc_hd__o21a_1
XANTENNA__2504__S _0220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1884_ VSS VDD _1358_ _1361_ _1026_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1909__A _1340_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1628__B _1173_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2505_ VSS VDD _0007_ _0443_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2436_ VDD VSS _1331_ _1320_ _1307_ core.ndc.row_out_n\[14\] VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__1644__A _1032_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1940__A2 _1395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2367_ VSS VDD _0377_ _0384_ _0383_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2298_ VSS VDD core.osr.next_result_w\[9\] _0321_ _0322_ VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_56_225 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2475__A core.pdc.row_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_72_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_21_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_21_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_247 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_269 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1729__A _1074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_en_bit_n[2] core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_30_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2221_ VSS VDD _0253_ core.cnb.result_out\[1\] _0254_ _0240_ VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_87_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2152_ VSS VDD _0194_ _0196_ _0195_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2083_ VDD VSS core.pdc.col_out_n\[21\] core.pdc.col_out\[21\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__2635__B1 _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2742__B _0637_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_21_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2985_ VSS VDD _0799_ _0875_ _0873_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1936_ VDD VSS _1284_ _1391_ _1393_ core.pdc.col_out\[0\] VSS VDD sky130_fd_sc_hd__a21o_1
X_1867_ VSS VDD _1349_ _1325_ core.ndc.row_bottotop_n\[5\] _1027_ core.pdc.row_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__o22a_2
X_1798_ VSS VDD _1272_ _1109_ _1298_ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk1\[27\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[27\] core.ndc.col_out_n\[27\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_88_158 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2419_ VDD VSS _0424_ core.osr.next_sample_count_w\[8\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_123_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_320 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_83_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_84_386 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_120_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_cgen_dlycontrol3_in[0] net19 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_79_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col_n[12] nmatrix_col_core_n_buffered\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_117 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1731__B _1188_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2562__B _0482_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2770_ VSS VDD _0656_ _0665_ _0666_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1721_ VDD VSS _1249_ _1246_ VSS VDD sky130_fd_sc_hd__inv_2
X_1652_ VDD VSS _1194_ _1193_ VSS VDD sky130_fd_sc_hd__inv_2
X_1583_ VDD VSS _1133_ _1132_ VSS VDD sky130_fd_sc_hd__inv_2
X_2204_ VSS VDD core.cnb.next_average_sum_w\[4\] _0238_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_3184_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0054_ net87 core.cnb.data_register_r\[4\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_2135_ VDD VSS core.cnb.average_counter_r\[3\] _0178_ core.cnb.average_counter_r\[4\]
+ _0179_ VSS VDD sky130_fd_sc_hd__a21o_1
X_2066_ VDD VSS _0139_ _1173_ core.pdc.col_out\[17\] _0089_ _1296_ _0140_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1831__A1 core.pdc.rowoff_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2968_ VSS VDD _0841_ _0852_ _0860_ _0859_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1919_ VSS VDD _1026_ _1029_ _1382_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_118_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2899_ VDD VSS _0792_ _0782_ _0775_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_134_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk2\[5\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[5\] core.ndc.rowon_bottotop_n\[5\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1551__B _1092_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_27_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk2\[0\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[0\] core.pdc.row_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_43_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_138_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2602__S _0438_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_197 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2066__B2 _1296_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2822_ VSS VDD _0714_ _0717_ _0716_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2753_ VDD VSS _0639_ _0649_ VSS VDD sky130_fd_sc_hd__buf_6
X_1704_ VSS VDD _1237_ core.ndc.col_out_n\[13\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1577__B1 _1082_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_69_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2684_ VDD VSS net39 core.osr.next_result_w\[6\] _0562_ _0586_ _0393_ VSS VDD sky130_fd_sc_hd__a22o_1
X_1635_ VDD VSS core.ndc.col_out\[7\] core.ndc.col_out_n\[7\] VSS VDD sky130_fd_sc_hd__inv_2
X_1566_ VSS VDD _1120_ _1110_ _1119_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1652__A _1193_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1497_ VSS VDD _1056_ _1057_ VSS VDD sky130_fd_sc_hd__clkbuf_4
X_3167_ VSS VDD net61 core.osr.next_result_w\[7\] net73 core.osr.result_r\[7\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_3098_ VSS VDD _0063_ _0980_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2118_ VSS VDD _0169_ _0168_ _0167_ _0166_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_120_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2049_ VSS VDD core.pdc.col_out_n\[14\] _0129_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_120_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_cgen_dlycontrol2_in[1] net30 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout57 VDD VSS net57 net58 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout68 VSS VDD net69 net68 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout79 VDD VSS net79 net80 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1562__A _1113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2377__B _0240_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_38_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_52 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2824__C core.cnb.pswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2599__A2 _0439_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_111 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1737__A _1074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1420_ VDD VSS core.osr.sample_count_r\[6\] core.osr.sample_count_r\[8\] core.osr.sample_count_r\[7\]
+ core.osr.sample_count_r\[4\] _0984_ VSS VDD sky130_fd_sc_hd__or4_1
XANTENNA__1472__A net15 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3021_ VSS VDD _0860_ _0909_ _0908_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2805_ VSS VDD _0645_ _0700_ _0642_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1647__A _1190_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2736_ VSS VDD _0630_ _0049_ _0632_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2667_ VSS VDD _0566_ _0570_ _0571_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1618_ VDD VSS _1164_ _1163_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1970__B1 _1045_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2598_ VSS VDD _1022_ _0509_ _0501_ _1328_ _0512_ _0461_ VSS VDD sky130_fd_sc_hd__o221a_1
XANTENNA__3190__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1549_ VSS VDD _1105_ _1056_ _1050_ VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_75_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_131_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1557__A _1085_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[8\].buf_p_rowonn_A core.pdc.rowon_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_215 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_92_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__3012__A _0799_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[9\].buf_n_rowonn_A core.ndc.rowon_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col[10] core.ndc.col_out\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2521_ VSS VDD _0452_ core.cnb.shift_register_r\[14\] _0219_ core.cnb.shift_register_r\[13\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_2452_ VDD VSS core.ndc.rowon_out_n\[12\] _0430_ VSS VDD sky130_fd_sc_hd__inv_2
X_2383_ VSS VDD core.osr.sample_count_r\[0\] core.osr.sample_count_r\[1\] _0396_ VSS
+ VDD sky130_fd_sc_hd__nor2_1
XANTENNA_cgen_dlycontrol1_in[2] net26 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_204 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xinput3 VSS VDD config_1_in[10] net3 VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1930__A core.pdc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3004_ VSS VDD _0892_ _0893_ _1117_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_281 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_101_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2480__B core.pdc.row_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2719_ VSS VDD _0517_ _0380_ _0617_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_126_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_120_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_87_521 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_42_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_92_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2581__A _0439_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1952_ VDD VSS _1406_ _1405_ VSS VDD sky130_fd_sc_hd__inv_2
X_1883_ VSS VDD _1360_ core.pdc.row_out_n\[14\] _1359_ VSS VDD sky130_fd_sc_hd__nor2_2
XANTENNA__1909__B core.pdc.rowoff_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2504_ VSS VDD _0443_ core.cnb.shift_register_r\[6\] _0220_ core.cnb.shift_register_r\[5\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_2435_ VSS VDD core.ndc.row_bottotop_n\[10\] _1318_ core.pdc.rowoff_out_n\[8\] _1369_
+ core.ndc.row_out_n\[13\] VSS VDD sky130_fd_sc_hd__o22a_1
X_2366_ VDD VSS _0383_ _0382_ VSS VDD sky130_fd_sc_hd__inv_2
X_2297_ VSS VDD _0252_ _0322_ core.cnb.result_out\[9\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_56_237 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk2\[5\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[5\] core.ndc.row_bottotop_n\[10\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1835__A net14 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_204 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_259 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk2\[13\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[13\] core.pdc.rowon_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1729__B _1243_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3101__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_en_bit_n[1] core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2220_ VDD VSS _0250_ _0249_ _0252_ _0253_ VSS VDD sky130_fd_sc_hd__a21o_1
Xpmat_sample_buf VSS VDD pmat_sample_switch_buffered net55 VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_23_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2151_ VDD VSS _0195_ _0177_ _0186_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_93_321 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2082_ VSS VDD _1284_ _0106_ _0148_ core.pdc.col_out_n\[21\] VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_93_376 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_387 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2635__A1 core.cnb.result_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2984_ VSS VDD _0874_ _0873_ _0784_ VSS VDD sky130_fd_sc_hd__or2_1
Xgenblk1\[0\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[0\] core.pdc.col_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1935_ VDD VSS _1393_ _1392_ VSS VDD sky130_fd_sc_hd__inv_2
X_1866_ VDD VSS _1349_ _1329_ VSS VDD sky130_fd_sc_hd__inv_2
X_1797_ VDD VSS core.ndc.col_out_n\[29\] core.ndc.col_out\[29\] VSS VDD sky130_fd_sc_hd__inv_2
X_2418_ VDD VSS _0423_ core.osr.is_last_sample _0422_ _0424_ VSS VDD sky130_fd_sc_hd__or3_1
XANTENNA__2486__A sample_nmatrix_cgen VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2349_ VDD VSS _0368_ core.osr.result_r\[15\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_84_332 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3124__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_99 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_79_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2396__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input33_A config_2_in[9] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[2\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[2\] core.ndc.row_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__3004__B _1117_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_368 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1720_ VDD VSS core.ndc.col_out\[15\] core.ndc.col_out_n\[15\] VSS VDD sky130_fd_sc_hd__inv_2
X_1651_ VSS VDD _1193_ _1192_ _1191_ _1077_ VSS VDD sky130_fd_sc_hd__o21a_2
XANTENNA__1475__A _1034_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1582_ VDD VSS _1113_ _1079_ _1051_ _1132_ VSS VDD sky130_fd_sc_hd__a21o_1
X_2203_ VSS VDD _0238_ _0237_ _0236_ _0209_ VSS VDD sky130_fd_sc_hd__and3_1
X_3183_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0053_ net86 core.cnb.data_register_r\[3\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_2134_ VSS VDD _0177_ _0178_ core.cnb.sampled_avg_control_r\[0\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_93_173 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2065_ VSS VDD _0065_ _1405_ _0140_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_139_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2967_ VSS VDD _0857_ _1076_ _0859_ _0858_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1918_ VSS VDD core.pdc.rowon_out_n\[10\] _1381_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2898_ VSS VDD _0789_ _0791_ _0790_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1849_ VDD VSS _1336_ _1026_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_118_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_76_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_138_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2066__A2 _1173_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_72_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2821_ VSS VDD _0471_ _0686_ _0716_ _0715_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2752_ VSS VDD _0648_ _0640_ _0647_ _0634_ VSS VDD sky130_fd_sc_hd__nand3b_1
X_1703_ VSS VDD _1237_ _1236_ _1234_ _1233_ VSS VDD sky130_fd_sc_hd__and3_1
X_2683_ VDD VSS _0581_ _0584_ _0585_ _0583_ VSS VDD sky130_fd_sc_hd__o21bai_1
X_1634_ VSS VDD _1179_ core.ndc.col_out_n\[7\] VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1565_ VSS VDD _1119_ _1118_ _1077_ _1112_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__1933__A _1057_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_405 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_58_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1496_ VSS VDD _1055_ _1056_ core.cnb.data_register_r\[3\] VSS VDD sky130_fd_sc_hd__nand2_1
X_3166_ VSS VDD net60 core.osr.next_result_w\[6\] net72 core.osr.result_r\[6\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_3097_ VSS VDD _0980_ core.osr.osr_mode_r\[1\] _0241_ net12 VSS VDD sky130_fd_sc_hd__mux2_1
X_2117_ VSS VDD _0077_ _0168_ _1235_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2048_ VSS VDD _0129_ _0128_ _0127_ _0123_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_120_48 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_cgen_dlycontrol2_in[0] net29 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xfanout58 VSS VDD net67 net58 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout69 VSS VDD net70 net69 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_13_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_129_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_129_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_64 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_70_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_79_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1472__B core.cnb.data_register_r\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3020_ VDD VSS _0908_ _0906_ _0907_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_95_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2804_ VSS VDD _0698_ _0699_ core.cnb.shift_register_r\[12\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_117_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2735_ VDD VSS _0632_ _0631_ VSS VDD sky130_fd_sc_hd__inv_2
X_2666_ VSS VDD _0567_ _0570_ _0569_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_2_1__f_clk_dig_dummy_A clknet_0_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1617_ VDD VSS _1163_ _1050_ _1162_ VSS VDD sky130_fd_sc_hd__or2_2
X_2597_ VSS VDD _0031_ _0511_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_115_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1548_ VSS VDD _1058_ _1104_ VSS VDD sky130_fd_sc_hd__clkbuf_4
X_1479_ VDD VSS _1039_ net15 VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_86_235 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3149_ VSS VDD net59 _0039_ net71 net49 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_54_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_131_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_360 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1573__A _1095_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_290 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[5\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[5\] core.pdc.col_out_n\[5\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2520_ VSS VDD _0014_ _0451_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2451_ VDD VSS _1328_ _1369_ _1365_ _0430_ _1331_ VSS VDD sky130_fd_sc_hd__a22o_1
X_2382_ VSS VDD _0395_ core.osr.next_sample_count_w\[0\] core.osr.sample_count_r\[0\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_dlycontrol1_in[1] net25 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_408 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput4 VSS VDD config_1_in[11] net4 VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1930__B _1040_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3003_ VSS VDD _0890_ _0892_ _0891_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_51_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_293 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2718_ VDD VSS _0616_ _0615_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_10_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2649_ VDD VSS _0394_ core.osr.next_result_w\[2\] _0542_ _0555_ net50 VSS VDD sky130_fd_sc_hd__a22o_1
XFILLER_86_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk2\[7\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[7\] core.ndc.row_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1568__A core.ndc.col_out_n\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2671__B _1002_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_129_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_76_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3180__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1951_ VSS VDD _1405_ _1403_ _1090_ _1404_ VSS VDD sky130_fd_sc_hd__a21bo_1
X_1882_ VSS VDD _1311_ _1349_ _1360_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2503_ VSS VDD _0006_ _0442_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2434_ VSS VDD _1325_ _1321_ core.pdc.rowoff_out_n\[8\] _1328_ core.ndc.row_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__o22a_1
X_2365_ VSS VDD core.osr.result_r\[16\] _0382_ core.osr.result_r\[17\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1689__B1 _1199_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1941__A _1396_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_503 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2296_ VSS VDD _0319_ _0271_ _0321_ _0320_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_2_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk1\[2\].buf_n_coln VDD VSS core.ndc.col_out_n\[2\] nmatrix_col_core_n_buffered\[2\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_52_488 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_137_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_137_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_216 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1570__B _1037_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_102_71 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_en_bit_n[0] core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3187__RESET_B net85 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1761__A _1072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2150_ VSS VDD _0192_ _0194_ _0190_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1480__B _1039_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2081_ VSS VDD _0075_ _0148_ _1284_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_93_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2983_ VSS VDD _0704_ _0873_ _0695_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_21_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1934_ VSS VDD _1390_ _1392_ _1069_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1865_ VDD VSS core.ndc.row_bottotop_n\[5\] _1348_ VSS VDD sky130_fd_sc_hd__inv_2
X_1796_ VDD VSS _1297_ _1296_ _1100_ _1091_ _1279_ core.ndc.col_out\[29\] VSS VDD
+ sky130_fd_sc_hd__a221o_2
XANTENNA__2571__A1 _0439_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2417_ VDD VSS _0423_ _0419_ core.osr.sample_count_r\[8\] VSS VDD sky130_fd_sc_hd__and2_1
X_2348_ VDD VSS core.osr.next_result_w\[14\] _0367_ VSS VDD sky130_fd_sc_hd__inv_2
X_2279_ VSS VDD core.osr.result_r\[8\] core.cnb.result_out\[8\] _0305_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_16_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[10] nmatrix_col_core_n_buffered\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1581__A _1039_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input26_A config_2_in[2] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_90_347 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1650_ VSS VDD _1077_ _1192_ _1132_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1581_ VSS VDD _1039_ _1131_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__2553__A1 core.cnb.result_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2202_ VSS VDD _0237_ _0235_ _0233_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_85_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3182_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0052_ net86 core.cnb.data_register_r\[2\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2133_ VSS VDD core.cnb.sampled_avg_control_r\[2\] _0176_ _0177_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_93_185 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2069__B1 _1075_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2064_ VDD VSS _0139_ _0125_ VSS VDD sky130_fd_sc_hd__inv_2
X_2966_ VSS VDD _0855_ _0858_ _0856_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1917_ VSS VDD _1381_ _1362_ core.ndc.rowoff_out_n\[5\] _1380_ VSS VDD sky130_fd_sc_hd__a21bo_1
X_2897_ VSS VDD _0786_ _0787_ _0790_ _1395_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1848_ VDD VSS core.pdc.row_out_n\[6\] _1335_ VSS VDD sky130_fd_sc_hd__inv_2
X_1779_ VDD VSS core.ndc.col_out_n\[25\] core.ndc.col_out\[25\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_76_119 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_94_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_138_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_rowoff_n[5] core.pdc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_92 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__3015__B _1312_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2820_ VSS VDD _0713_ _0715_ VSS VDD sky130_fd_sc_hd__clkinvlp_2
XFILLER_129_143 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2751_ VSS VDD _0643_ _0646_ _0647_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2682_ VSS VDD core.osr.next_result_w\[8\] _0540_ _0584_ _0528_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1702_ VSS VDD _1149_ _1236_ _1235_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1577__A2 _1128_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1486__A _1045_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1633_ VSS VDD _1179_ _1178_ _1174_ _1168_ VSS VDD sky130_fd_sc_hd__and3_1
X_1564_ VSS VDD _1116_ _1118_ _1117_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1495_ VDD VSS _1055_ core.cnb.data_register_r\[4\] VSS VDD sky130_fd_sc_hd__buf_4
XANTENNA__3114__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3165_ VSS VDD net60 core.osr.next_result_w\[5\] net72 core.osr.result_r\[5\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_66_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3096_ VSS VDD _0062_ _0979_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2116_ VSS VDD _1406_ _0167_ _1188_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2047_ VSS VDD _1413_ _0128_ _1235_ VSS VDD sky130_fd_sc_hd__nand2_1
Xfanout59 VDD VSS net59 net61 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2949_ VSS VDD _0839_ _0482_ _0841_ _0840_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_129_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2004__B _1284_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk1\[17\].buf_n_coln_A core.ndc.col_out_n\[17\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout76_A net82 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_32 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_110_60 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[1\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[1\] core.ndc.rowon_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_70_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3137__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[7\].buf_n_coln VDD VSS core.ndc.col_out_n\[7\] nmatrix_col_core_n_buffered\[7\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_2803_ VDD VSS _0698_ core.cnb.shift_register_r\[13\] VSS VDD sky130_fd_sc_hd__inv_2
X_2734_ VDD VSS _0393_ core.cnb.result_out\[11\] _0562_ _0631_ net44 VSS VDD sky130_fd_sc_hd__a22o_1
X_2665_ VSS VDD core.osr.next_result_w\[8\] _0569_ _0568_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2596_ VSS VDD _0511_ core.cnb.result_out\[9\] _0480_ _0510_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1616_ VDD VSS _1162_ _1036_ _1134_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_115_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1547_ VSS VDD _1078_ _1103_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1478_ VSS VDD _1031_ _1038_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3148_ VSS VDD net56 _0038_ net68 net48 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3079_ VSS VDD _0965_ _0955_ _0964_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_24_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_108_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1748__B _1173_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2450_ VSS VDD _1378_ core.ndc.rowon_out_n\[11\] _1370_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2381_ VDD VSS _0395_ _0394_ VSS VDD sky130_fd_sc_hd__buf_4
XANTENNA_cgen_dlycontrol1_in[0] net18 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput5 VSS VDD config_1_in[12] net5 VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3002_ VSS VDD _0847_ _0891_ _0888_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_91_261 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2534__S net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2717_ VDD VSS core.osr.next_result_w\[10\] net43 _0393_ _0615_ _0562_ VSS VDD sky130_fd_sc_hd__a22o_1
X_2648_ VSS VDD _0554_ _0516_ _0520_ VSS VDD sky130_fd_sc_hd__or2_1
X_2579_ VDD VSS _0027_ _0496_ _0497_ _0461_ core.cnb.result_out\[5\] VSS VDD sky130_fd_sc_hd__o2bb2a_1
XFILLER_47_409 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_453 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_136 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1950_ VSS VDD _1400_ _1404_ _1086_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1881_ VSS VDD _1336_ _1358_ _1359_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2502_ VSS VDD _0442_ core.cnb.shift_register_r\[5\] _0203_ core.cnb.shift_register_r\[4\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__2583__C1 _0439_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2433_ VDD VSS core.ndc.row_out_n\[11\] _0427_ VSS VDD sky130_fd_sc_hd__inv_2
X_2364_ VDD VSS core.osr.result_r\[16\] _0377_ core.osr.result_r\[17\] _0381_ VSS
+ VDD sky130_fd_sc_hd__a21o_1
XFILLER_110_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2295_ VSS VDD _0318_ _0320_ _0317_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_84_515 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2491__C _1040_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3095__S _0241_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_342 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_127_91 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2080_ VDD VSS core.pdc.col_out_n\[20\] core.pdc.col_out\[20\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_93_367 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2096__B2 _1102_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1489__A _1037_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2982_ VSS VDD _0055_ _0757_ _0872_ _0871_ _1114_ _0688_ VSS VDD sky130_fd_sc_hd__a32o_1
X_1933_ VDD VSS _1089_ _1390_ _1057_ _1391_ VSS VDD sky130_fd_sc_hd__or3_1
X_1864_ VSS VDD _1308_ _1318_ _1348_ VSS VDD sky130_fd_sc_hd__nor2_1
Xinput30 VDD VSS net30 config_2_in[6] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_1795_ VSS VDD _1272_ _1143_ _1297_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2416_ VSS VDD core.osr.sample_count_r\[8\] _0419_ _0422_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2347_ VSS VDD _0365_ _0240_ _0367_ _0366_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2278_ VSS VDD _0304_ core.osr.next_result_w\[7\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_16_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_79_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__3170__CLK net61 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2693__A _0395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input19_A config_2_in[10] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1580_ VDD VSS core.ndc.col_out_n\[4\] core.ndc.col_out\[4\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2002__A1 _1082_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2201_ VSS VDD _0233_ _0236_ _0235_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3181_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0051_ net86 core.cnb.data_register_r\[1\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_4
X_2132_ VDD VSS _0176_ core.cnb.sampled_avg_control_r\[1\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2069__A1 _1126_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2069__B2 _0115_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2063_ VDD VSS core.pdc.col_out_n\[16\] core.pdc.col_out\[16\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__2108__A _1131_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2965_ VDD VSS _0855_ _0831_ _0856_ _0857_ VSS VDD sky130_fd_sc_hd__a21o_1
X_1916_ VSS VDD _1372_ _1380_ _1331_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2896_ VSS VDD _0788_ _0789_ _1076_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1847_ VDD VSS _1331_ _1320_ _1334_ _1335_ VSS VDD sky130_fd_sc_hd__a21o_1
X_1778_ VSS VDD core.ndc.col_out\[25\] _1157_ _1284_ _1285_ _1287_ VSS VDD sky130_fd_sc_hd__a211o_2
XANTENNA_genblk2\[5\].buf_p_rown_A core.ndc.row_bottotop_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_138_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1576__B _1057_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_84_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1767__A _1032_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2750_ VSS VDD _0646_ _0644_ _0645_ VSS VDD sky130_fd_sc_hd__nand2_2
X_2681_ VSS VDD _0356_ _0582_ _0583_ _0517_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1701_ VDD VSS _1235_ net15 VSS VDD sky130_fd_sc_hd__buf_2
X_1632_ VSS VDD _1176_ _1178_ _1177_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__3171__RESET_B net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1563_ VDD VSS _1117_ core.cnb.data_register_r\[7\] VSS VDD sky130_fd_sc_hd__buf_2
X_1494_ VSS VDD _1041_ _1054_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__2110__B _1177_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3164_ VSS VDD net62 core.osr.next_result_w\[4\] net74 core.osr.result_r\[4\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_3095_ VSS VDD _0979_ core.osr.osr_mode_r\[0\] _0241_ net11 VSS VDD sky130_fd_sc_hd__mux2_1
X_2115_ VSS VDD _1398_ _0166_ _1096_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2046_ VDD VSS _0126_ _0127_ VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1677__A _1216_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2948_ VDD VSS _0840_ _0791_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_129_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_135_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2879_ VSS VDD _0771_ _0773_ _0772_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2020__B _1093_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_85_462 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_85_495 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_110_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_70_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_79_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2802_ VSS VDD _0684_ _0696_ _0697_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2733_ VSS VDD _0628_ _0630_ _0629_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2105__B _1092_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2664_ VSS VDD _1001_ _0568_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2595_ VSS VDD _0510_ _0508_ _0509_ VSS VDD sky130_fd_sc_hd__or2_1
X_1615_ VSS VDD _1160_ _1161_ _1051_ VSS VDD sky130_fd_sc_hd__nor2_2
Xgenblk2\[6\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[6\] core.pdc.rowon_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA_cgen_enable_dlycontrol_in net24 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1546_ VDD VSS _1102_ _1101_ VSS VDD sky130_fd_sc_hd__buf_2
X_1477_ VDD VSS _1037_ _1036_ VSS VDD sky130_fd_sc_hd__inv_2
X_3147_ VSS VDD net56 _0037_ net68 net47 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3078_ VSS VDD _0957_ _0964_ _0963_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2435__B2 core.ndc.row_bottotop_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2435__A1 core.pdc.rowoff_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2029_ VSS VDD _0084_ _0114_ _1155_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_genblk2\[15\].buf_p_rowonn_A core.pdc.rowon_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_88 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3104__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_81_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2380_ VSS VDD _0393_ _0394_ VSS VDD sky130_fd_sc_hd__clkbuf_2
Xinput6 VSS VDD config_1_in[13] net6 VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3001_ VSS VDD _0795_ _0890_ _0889_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_229 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_101_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2716_ VSS VDD _0612_ _0047_ _0614_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2647_ VDD VSS _1000_ core.osr.next_result_w\[10\] _0552_ _0553_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__1674__B _1213_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2578_ VDD VSS _1065_ _0489_ _0480_ _0497_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_1529_ VDD VSS _1087_ _1044_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__3127__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_67 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_89 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_row_n[1] nmatrix_row_core_n_buffered\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_76_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_112 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1880_ VSS VDD _1317_ _1358_ _1029_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1775__A _1126_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2501_ VSS VDD _0005_ _0441_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2432_ VSS VDD _1322_ _0427_ _1330_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2363_ VDD VSS core.osr.next_result_w\[16\] _0380_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1689__A2 _1206_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2294_ VSS VDD _0319_ _0317_ _0318_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_112_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_137_37 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_295 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_15_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1595__A _1045_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2096__A2 _1275_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_262 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_295 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2981_ VSS VDD _0863_ _0802_ _0872_ _0870_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1932_ VDD VSS _1390_ _1389_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_1863_ VDD VSS core.pdc.row_out_n\[9\] _1347_ VSS VDD sky130_fd_sc_hd__inv_2
Xinput31 VDD VSS net31 config_2_in[7] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 VDD VSS net20 config_2_in[11] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_1794_ VDD VSS _1296_ _1095_ VSS VDD sky130_fd_sc_hd__buf_2
X_2415_ VDD VSS core.osr.next_sample_count_w\[7\] _0421_ VSS VDD sky130_fd_sc_hd__inv_2
X_2346_ VSS VDD _0353_ core.osr.result_r\[14\] _0366_ _0358_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2277_ VSS VDD core.cnb.result_out\[7\] _0271_ _0303_ _0304_ VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_12_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_316 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_113_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_73_76 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2200_ VDD VSS _0235_ core.cnb.average_sum_r\[4\] VSS VDD sky130_fd_sc_hd__inv_2
X_3180_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0050_ net86 core.cnb.data_register_r\[0\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_4
X_2131_ VDD VSS core.cnb.data_register_r\[2\] core.cnb.pswitch_out\[2\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2062_ VSS VDD _1075_ _0135_ _0094_ _1064_ core.pdc.col_out_n\[16\] _0138_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_75_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2108__B _0091_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2964_ VSS VDD _0847_ _0856_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1915_ VSS VDD core.ndc.rowoff_out_n\[5\] core.ndc.row_bottotop_n\[5\] core.ndc.rowon_bottotop_n\[5\]
+ VSS VDD sky130_fd_sc_hd__nand2_2
X_2895_ VSS VDD _0786_ _0788_ _0787_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1846_ VSS VDD _1333_ _1316_ _1334_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1777_ VDD VSS _1287_ _1286_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_89_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1504__A1 _1035_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2329_ VSS VDD _0351_ _0317_ _0307_ _0350_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_66_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1873__A _1353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1592__B _1112_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_87 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input31_A config_2_in[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_84_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_72_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2680_ VSS VDD core.osr.next_result_w\[10\] _0582_ _0568_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1700_ VSS VDD _1234_ _1034_ _1204_ VSS VDD sky130_fd_sc_hd__or2_1
X_1631_ VDD VSS _1177_ _1072_ VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1783__A _1131_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1562_ VSS VDD _1113_ _1115_ _1116_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1493_ VSS VDD _1052_ _1053_ VSS VDD sky130_fd_sc_hd__clkbuf_4
X_3163_ VSS VDD net63 core.osr.next_result_w\[3\] net74 core.osr.result_r\[3\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__3140__RESET_B net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2114_ VDD VSS core.pdc.col_out_n\[28\] core.pdc.col_out\[28\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_3094_ VSS VDD _0977_ _0061_ _0978_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_81_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2045_ VSS VDD _1227_ _0125_ _0126_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_63_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2947_ VDD VSS _0475_ _0837_ _0838_ _0839_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_129_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2878_ VSS VDD _0772_ _0471_ _0760_ _0770_ VSS VDD sky130_fd_sc_hd__nand3b_1
XANTENNA__1973__B2 _1296_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1973__A1 _1121_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_135_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1829_ VSS VDD _1022_ _1319_ _1320_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_79_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_135_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_63_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3183__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2801_ VSS VDD _0693_ _0696_ _0695_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2732_ VDD VSS _0530_ _0363_ _1018_ _0629_ VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__1955__B2 _1296_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2663_ VSS VDD core.osr.next_result_w\[10\] _0567_ _0535_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2594_ VSS VDD _1303_ _0503_ _0509_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1614_ VSS VDD _1058_ _1066_ _1160_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1545_ VSS VDD _1032_ _1101_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__2121__B _1096_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1476_ VSS VDD _1036_ core.cnb.data_register_r\[3\] core.cnb.data_register_r\[4\]
+ VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_86_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3146_ VSS VDD net56 _0036_ net68 net46 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_54_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3077_ VSS VDD _0948_ _0960_ _0962_ _0963_ VSS VDD sky130_fd_sc_hd__o21a_1
X_2028_ VSS VDD _1136_ _1228_ _0113_ _1394_ VSS VDD sky130_fd_sc_hd__o21ai_2
XANTENNA__1688__A _1074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2791__B core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1643__B1 _1186_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A net82 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_81_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_81_76 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk1\[13\].buf_n_coln_A core.ndc.col_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_107 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2222__A _0254_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1780__B _1284_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput7 VSS VDD config_1_in[14] net7 VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3000_ VDD VSS _0889_ _0888_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2116__B _1188_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[13\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[13\] core.pdc.row_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2715_ VDD VSS _0614_ _0613_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2132__A core.cnb.sampled_avg_control_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2646_ VSS VDD _0550_ _0552_ _0551_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2577_ VSS VDD _0493_ _0496_ _1114_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1690__B _1093_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1528_ VSS VDD _1079_ _1085_ _1086_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1459_ VDD VSS core.cnb.data_register_r\[10\] _1022_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_27_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3129_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[2\] net91
+ core.cnb.average_sum_r\[2\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_55_455 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_160 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2042__A _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_row_n[0] nmatrix_row_core_n_buffered\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2032__A0 _1199_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2500_ VSS VDD _0441_ core.cnb.shift_register_r\[4\] _0220_ core.cnb.shift_register_r\[3\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__2583__B2 _1117_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2431_ VSS VDD core.ndc.row_bottotop_n\[10\] _1321_ _1311_ _1027_ core.ndc.row_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__o22a_1
XANTENNA__1791__A _1272_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2362_ VSS VDD _0378_ _0241_ _0380_ _0379_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2293_ VSS VDD _0311_ _0318_ _0306_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_56_208 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_sample_buf_n_A core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1966__A core.pdc.col_out\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2629_ VDD VSS _0537_ _1011_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_102_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2037__A _0098_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[10\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[10\] core.ndc.row_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1595__B _1079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_119 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1525__C1 _1082_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[15\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[15\] core.ndc.rowon_out_n\[15\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_46_230 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2980_ VDD VSS _0802_ _0863_ _0870_ _0871_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__1786__A _1106_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1931_ VSS VDD _1388_ _1389_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1862_ VDD VSS _1347_ _1344_ _1346_ VSS VDD sky130_fd_sc_hd__or2_2
Xinput21 VDD VSS net21 config_2_in[12] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 VSS VDD net10 config_1_in[2] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2005__B1 _1035_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1793_ VDD VSS core.ndc.col_out_n\[28\] core.ndc.col_out\[28\] VSS VDD sky130_fd_sc_hd__inv_2
Xinput32 VDD VSS net32 config_2_in[8] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2414_ VSS VDD _1021_ _0420_ _0419_ _0421_ VSS VDD sky130_fd_sc_hd__or3b_1
XANTENNA__3117__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2345_ VSS VDD _0359_ _0365_ _0364_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2276_ VSS VDD _0302_ _0255_ _0303_ _0301_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_84_369 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_506 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_328 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_73_88 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_92 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_98_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[14\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[14\] core.pdc.col_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2230__A _0255_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3045__B _1114_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2130_ VDD VSS core.pdc.col_out\[31\] core.pdc.col_out_n\[31\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_14_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2061_ VSS VDD _1391_ _0138_ _1093_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2963_ VSS VDD _0855_ _0818_ _0745_ _0854_ VSS VDD sky130_fd_sc_hd__and3_1
X_1914_ VSS VDD _1336_ _1366_ core.pdc.rowon_out_n\[9\] core.ndc.rowon_bottotop_n\[5\]
+ VSS VDD sky130_fd_sc_hd__a21oi_2
X_2894_ VSS VDD _0787_ _0783_ _0472_ _0785_ VSS VDD sky130_fd_sc_hd__nand3b_1
X_1845_ VSS VDD _1332_ _1333_ _1300_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1776_ VSS VDD _1286_ _1033_ _1119_ VSS VDD sky130_fd_sc_hd__or2_1
X_2328_ VSS VDD _0332_ _0344_ _0350_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_84_111 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2259_ VSS VDD _0288_ _0287_ _0240_ _0280_ VSS VDD sky130_fd_sc_hd__o21a_2
XFILLER_43_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2985__A _0799_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_99 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_88_494 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input24_A config_2_in[15] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1630_ VDD VSS _1176_ _1175_ VSS VDD sky130_fd_sc_hd__inv_2
X_1561_ VSS VDD _1114_ _1037_ _1115_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1492_ VSS VDD _1051_ _1052_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3162_ VSS VDD net63 core.osr.next_result_w\[2\] net75 core.osr.result_r\[2\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2113_ VSS VDD core.pdc.col_out_n\[28\] _0165_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_3093_ VSS VDD _0758_ _0978_ _1309_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__3180__RESET_B net86 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2044_ VSS VDD _1161_ _1403_ _0124_ _0125_ VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_50_501 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2946_ VSS VDD _0475_ _0835_ _0838_ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk1\[11\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[11\] core.ndc.col_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2877_ VSS VDD _0761_ _0771_ _0770_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_135_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1828_ VDD VSS _1319_ _1028_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1974__A core.pdc.col_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_135_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1759_ VDD VSS core.ndc.col_out_n\[22\] core.ndc.col_out\[22\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col[9] core.ndc.col_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2029__B _1155_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[1\].buf_p_rown_A core.pdc.row_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2045__A _1227_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_110_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_144 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_63_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2881__C _0482_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2800_ VSS VDD _0640_ _0682_ _0695_ _0694_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2731_ VSS VDD _0623_ _0628_ _0627_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1794__A _1095_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1955__A2 _1279_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_117_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2662_ VDD VSS _1008_ _0356_ _0524_ _0566_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_1613_ VDD VSS core.ndc.col_out_n\[6\] core.ndc.col_out\[6\] VSS VDD sky130_fd_sc_hd__inv_2
X_2593_ VSS VDD _0507_ _0502_ _0508_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_132_119 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1544_ VDD VSS _1100_ _1099_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_5_84 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1475_ VDD VSS _1035_ _1034_ VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__2668__B1 _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3145_ VSS VDD net56 _0035_ net68 net45 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3076_ VSS VDD _0962_ _0961_ _0833_ _0918_ _0507_ VSS VDD sky130_fd_sc_hd__a211o_1
X_2027_ VDD VSS core.pdc.col_out_n\[11\] core.pdc.col_out\[11\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_50_331 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1643__A1 _1113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2929_ VDD VSS _0821_ _0818_ VSS VDD sky130_fd_sc_hd__inv_2
Xgenblk2\[15\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[15\] core.ndc.row_out_n\[15\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_108_116 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_40_37 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_123_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_35 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_105_74 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_45_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_128 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_81_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_114_119 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_122_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput8 VSS VDD config_1_in[15] net8 VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_51_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2714_ VDD VSS core.osr.next_result_w\[9\] net42 _1020_ _0613_ _0562_ VSS VDD sky130_fd_sc_hd__a22o_1
X_2645_ VDD VSS _1001_ core.osr.next_result_w\[6\] _1009_ _0551_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_10_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2576_ VSS VDD _0026_ _0495_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2889__B1 _0482_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1527_ VDD VSS _1085_ _1081_ VSS VDD sky130_fd_sc_hd__buf_2
X_1458_ VSS VDD _1021_ core.osr.is_last_sample VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3128_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[1\] net90
+ core.cnb.average_sum_r\[1\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_27_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_423 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3059_ VSS VDD _0946_ _0507_ _0945_ VSS VDD sky130_fd_sc_hd__or2_1
Xgenblk2\[2\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[2\] core.pdc.rowon_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_51_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2042__B _1279_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3173__CLK net61 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[19\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[19\] core.pdc.col_out_n\[19\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_18_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_412 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_434 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_41_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2583__A2 _1067_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2430_ VDD VSS _0426_ core.ndc.row_bottotop_n\[10\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1791__B _1175_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2361_ VSS VDD _0377_ _0379_ core.osr.result_r\[16\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2292_ VSS VDD _0314_ _0316_ _0317_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2099__A1 _0081_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2099__B2 _1096_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[21\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[21\] core.pdc.col_out_n\[21\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_52_437 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2628_ VSS VDD core.osr.next_result_w\[6\] _0536_ _0535_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2559_ VSS VDD _0023_ _0481_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_46_36 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_102_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_337 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_286 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1930_ VSS VDD core.pdc.rowon_out_n\[0\] _1388_ _1040_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1861_ VDD VSS _1346_ _1345_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1786__B _1188_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput22 VDD VSS net22 config_2_in[13] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_90 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput11 VSS VDD net11 config_1_in[3] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2005__B2 _0072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2005__A1 _1126_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[16\].buf_n_coln VDD VSS core.ndc.col_out_n\[16\] nmatrix_col_core_n_buffered\[16\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_1792_ VDD VSS _1295_ _1125_ _1240_ _1294_ _1279_ core.ndc.col_out\[28\] VSS VDD
+ sky130_fd_sc_hd__a221o_2
Xinput33 VDD VSS net33 config_2_in[9] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_2413_ VSS VDD _0417_ _0420_ _1013_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_88_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2344_ VDD VSS _0364_ core.osr.result_r\[14\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_96_120 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2275_ VSS VDD _0302_ _0300_ _0290_ _0294_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_92_392 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_32_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_57_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_518 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_57_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_73_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1994__A0 _1202_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_98_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2060_ VDD VSS core.pdc.col_out_n\[15\] core.pdc.col_out\[15\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1797__A core.ndc.col_out\[29\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2962_ VSS VDD _0854_ _0737_ _0734_ _0853_ VSS VDD sky130_fd_sc_hd__and3_1
X_1913_ VSS VDD core.pdc.rowon_out_n\[8\] _1379_ core.ndc.rowon_out_n\[15\] VSS VDD
+ sky130_fd_sc_hd__nand2_2
X_2893_ VSS VDD _0784_ _0786_ _0785_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_8_62 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1844_ VSS VDD _1303_ _1326_ _1332_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1775_ VSS VDD _1126_ _1231_ _1285_ VSS VDD sky130_fd_sc_hd__nor2_1
Xnmat nmatrix_row_core_n_buffered\[0\] nmatrix_row_core_n_buffered\[1\] nmatrix_row_core_n_buffered\[2\]
+ nmatrix_row_core_n_buffered\[3\] nmatrix_row_core_n_buffered\[4\] nmatrix_row_core_n_buffered\[5\]
+ nmatrix_row_core_n_buffered\[6\] nmatrix_row_core_n_buffered\[7\] nmatrix_row_core_n_buffered\[8\]
+ nmatrix_row_core_n_buffered\[9\] nmatrix_row_core_n_buffered\[10\] nmatrix_row_core_n_buffered\[11\]
+ nmatrix_row_core_n_buffered\[12\] nmatrix_row_core_n_buffered\[13\] nmatrix_row_core_n_buffered\[14\]
+ nmatrix_row_core_n_buffered\[15\] nmatrix_rowon_core_n_buffered\[0\] nmatrix_rowon_core_n_buffered\[1\]
+ nmatrix_rowon_core_n_buffered\[2\] nmatrix_rowon_core_n_buffered\[3\] nmatrix_rowon_core_n_buffered\[4\]
+ nmatrix_rowon_core_n_buffered\[5\] nmatrix_rowon_core_n_buffered\[6\] nmatrix_rowon_core_n_buffered\[7\]
+ nmatrix_rowon_core_n_buffered\[8\] nmatrix_rowon_core_n_buffered\[9\] nmatrix_rowon_core_n_buffered\[10\]
+ nmatrix_rowon_core_n_buffered\[11\] nmatrix_rowon_core_n_buffered\[12\] nmatrix_rowon_core_n_buffered\[13\]
+ nmatrix_rowon_core_n_buffered\[14\] nmatrix_rowon_core_n_buffered\[15\] core.ndc.rowoff_out_n\[0\]
+ core.ndc.rowoff_out_n\[1\] core.ndc.rowoff_out_n\[2\] core.ndc.rowoff_out_n\[3\]
+ core.ndc.rowoff_out_n\[4\] core.ndc.rowoff_out_n\[5\] core.ndc.rowoff_out_n\[6\]
+ core.ndc.rowoff_out_n\[7\] core.ndc.rowoff_out_n\[8\] core.ndc.rowoff_out_n\[9\]
+ core.ndc.rowoff_out_n\[10\] core.ndc.rowoff_out_n\[11\] core.ndc.rowoff_out_n\[12\]
+ core.ndc.rowoff_out_n\[13\] core.ndc.rowoff_out_n\[14\] core.ndc.rowoff_out_n\[15\]
+ vcm/vcm sample_nmatrix_cgen _0001_ nmatrix_col_core_n_buffered\[31\] nmatrix_col_core_n_buffered\[30\]
+ nmatrix_col_core_n_buffered\[29\] nmatrix_col_core_n_buffered\[28\] nmatrix_col_core_n_buffered\[27\]
+ nmatrix_col_core_n_buffered\[26\] nmatrix_col_core_n_buffered\[25\] nmatrix_col_core_n_buffered\[24\]
+ nmatrix_col_core_n_buffered\[23\] nmatrix_col_core_n_buffered\[22\] nmatrix_col_core_n_buffered\[21\]
+ nmatrix_col_core_n_buffered\[20\] nmatrix_col_core_n_buffered\[19\] nmatrix_col_core_n_buffered\[18\]
+ nmatrix_col_core_n_buffered\[17\] nmatrix_col_core_n_buffered\[16\] nmatrix_col_core_n_buffered\[15\]
+ nmatrix_col_core_n_buffered\[14\] nmatrix_col_core_n_buffered\[13\] nmatrix_col_core_n_buffered\[12\]
+ nmatrix_col_core_n_buffered\[11\] nmatrix_col_core_n_buffered\[10\] nmatrix_col_core_n_buffered\[9\]
+ nmatrix_col_core_n_buffered\[8\] nmatrix_col_core_n_buffered\[7\] nmatrix_col_core_n_buffered\[6\]
+ nmatrix_col_core_n_buffered\[5\] nmatrix_col_core_n_buffered\[4\] nmatrix_col_core_n_buffered\[3\]
+ nmatrix_col_core_n_buffered\[2\] nmatrix_col_core_n_buffered\[1\] nmatrix_col_core_n_buffered\[0\]
+ core.cnb.pswitch_out\[2\] core.cnb.pswitch_out\[1\] core.cnb.pswitch_out\[0\] net96
+ nmat_sample_switch_buffered nmat_sample_switch_n_buffered inn_analog core.ndc.col_out\[0\]
+ core.ndc.col_out\[1\] core.ndc.col_out\[2\] core.ndc.col_out\[3\] core.ndc.col_out\[4\]
+ core.ndc.col_out\[5\] core.ndc.col_out\[6\] core.ndc.col_out\[7\] core.ndc.col_out\[8\]
+ core.ndc.col_out\[9\] core.ndc.col_out\[10\] core.ndc.col_out\[11\] core.ndc.col_out\[12\]
+ core.ndc.col_out\[13\] core.ndc.col_out\[14\] core.ndc.col_out\[15\] core.ndc.col_out\[16\]
+ core.ndc.col_out\[17\] core.ndc.col_out\[18\] core.ndc.col_out\[19\] core.ndc.col_out\[20\]
+ core.ndc.col_out\[21\] core.ndc.col_out\[22\] core.ndc.col_out\[23\] core.ndc.col_out\[24\]
+ core.ndc.col_out\[25\] core.ndc.col_out\[26\] core.ndc.col_out\[27\] core.ndc.col_out\[28\]
+ core.ndc.col_out\[29\] core.ndc.col_out\[30\] core.ndc.col_out\[31\] ctop_nmatrix_analog
+ VSS VDD adc_array_matrix_12bit
X_2327_ VSS VDD core.osr.next_result_w\[11\] _0349_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2258_ VSS VDD _0285_ _0271_ _0287_ _0286_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_84_123 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_145 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2189_ VDD VSS _0226_ core.cnb.average_sum_r\[2\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1500__A _1057_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1976__A0 _1197_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_108_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_input17_A config_1_in[9] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_99 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2506__A _0208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3107__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1719__B1 _1075_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1560_ VDD VSS _1114_ _1044_ VSS VDD sky130_fd_sc_hd__buf_2
Xclkbuf_2_2__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_2__leaf_clk_dig_dummy
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
X_1491_ VSS VDD _1050_ _1051_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_3161_ VSS VDD net62 core.osr.next_result_w\[1\] net74 core.osr.result_r\[1\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2112_ VSS VDD _0165_ _0164_ _0163_ _0162_ VSS VDD sky130_fd_sc_hd__and3_1
X_3092_ VSS VDD _0976_ _0977_ _0689_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_54_329 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2043_ VSS VDD _1403_ _0124_ _1163_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_50_513 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2945_ VSS VDD _0831_ _0837_ _0836_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1958__B1 _1047_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2876_ VSS VDD _0769_ _0768_ _0764_ _0770_ VSS VDD sky130_fd_sc_hd__nor3_1
X_1827_ VSS VDD _1317_ _1318_ core.cnb.data_register_r\[10\] VSS VDD sky130_fd_sc_hd__nand2_1
X_1758_ VDD VSS _1273_ _1125_ _1217_ _1121_ _1193_ core.ndc.col_out\[22\] VSS VDD
+ sky130_fd_sc_hd__a221o_2
X_1689_ VSS VDD _1206_ _1103_ _1225_ _1199_ VSS VDD sky130_fd_sc_hd__a21oi_2
XANTENNA_nmat_col[8] core.ndc.col_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input9_A config_1_in[1] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2045__B _0125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2996__A _1113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_435 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[26\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[26\] core.pdc.col_out_n\[26\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2730_ VSS VDD _0530_ _0626_ _0627_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2661_ VSS VDD core.osr.next_result_w\[6\] _0540_ _0565_ _0528_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1612_ VDD VSS _1154_ core.ndc.col_out\[6\] _1152_ _1159_ _1155_ _1157_ VSS VDD sky130_fd_sc_hd__a221o_4
XFILLER_5_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2592_ VDD VSS _0507_ core.cnb.data_register_r\[9\] VSS VDD sky130_fd_sc_hd__inv_2
X_1543_ VSS VDD _1099_ _1067_ _1054_ _1098_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_5_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1474_ VDD VSS _1034_ _1033_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_39_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3144_ VSS VDD net56 _0034_ net68 net38 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3075_ VDD VSS _0833_ _0831_ _0918_ _0961_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_54_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2026_ VSS VDD _1064_ _0111_ _0110_ _1224_ core.pdc.col_out_n\[11\] _0112_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_90_490 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1985__A _0081_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2928_ VSS VDD _0819_ _0809_ _0806_ _0820_ VSS VDD sky130_fd_sc_hd__nor3_1
XANTENNA_genblk1\[9\].buf_n_coln_A core.ndc.col_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2859_ VSS VDD core.cnb.pswitch_out\[0\] _0753_ _0754_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_108_128 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_116_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_105_86 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_192 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2056__A _1242_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_dig_dummy_A clknet_0_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_122_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_genblk2\[14\].buf_p_rown_A core.pdc.row_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput9 VSS VDD net9 config_1_in[1] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_49_487 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2713_ VSS VDD _0610_ _0540_ _0612_ _0611_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2644_ VSS VDD core.osr.next_result_w\[8\] _0550_ _1002_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_65_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2575_ VSS VDD _0495_ core.cnb.result_out\[4\] _0480_ _0494_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1526_ VDD VSS _1084_ _1083_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2889__B2 _0758_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1457_ VDD VSS _1021_ _1020_ VSS VDD sky130_fd_sc_hd__inv_2
X_3127_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[0\] net90
+ core.cnb.average_sum_r\[0\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_27_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[23\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[23\] core.ndc.col_out_n\[23\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_55_479 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3058_ VSS VDD _0945_ _0799_ _0693_ _0472_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2009_ VDD VSS _0099_ _0100_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_136_7 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_116_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1552__A1 _1091_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1552__B2 _1102_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_479 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2360_ VSS VDD _0378_ core.osr.result_r\[16\] _0377_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1543__A1 _1067_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2291_ VDD VSS _0316_ _0315_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2099__A2 _1173_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2627_ VSS VDD _1002_ _0535_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2558_ VSS VDD _0481_ core.cnb.result_out\[1\] _0480_ _0479_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2489_ VSS VDD net64 _0435_ core.osr.data_valid_r VSS VDD sky130_fd_sc_hd__nand2_1
X_1509_ VSS VDD _1067_ _1046_ _1066_ VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__2318__B core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3140__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2988__B _1113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1525__A1 _1076_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_349 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1860_ VDD VSS core.cnb.data_register_r\[8\] _1304_ core.cnb.data_register_r\[11\]
+ net14 _1345_ VSS VDD sky130_fd_sc_hd__or4_1
Xinput12 VSS VDD net12 config_1_in[4] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1791_ VSS VDD _1272_ _1175_ _1295_ VSS VDD sky130_fd_sc_hd__nor2_1
Xinput23 VDD VSS net23 config_2_in[14] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 VSS VDD net34 rst_n VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2412_ VSS VDD _1013_ _0417_ _0419_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2343_ VDD VSS core.osr.next_result_w\[13\] _0363_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__3103__RESET_B net85 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_132 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2274_ VDD VSS _0290_ _0294_ _0300_ _0301_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_78_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1989_ VSS VDD _0086_ _0085_ _0082_ _0080_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_57_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_69_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_87_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_87_176 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_113_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_24 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1691__B1 _1035_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2064__A _0125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1994__A1 _1242_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_136 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[1\].buf_p_rowonn_A core.pdc.rowon_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_genblk2\[2\].buf_n_rowonn_A core.ndc.rowon_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3186__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1682__B1 _1137_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2961_ VDD VSS _0853_ _0742_ VSS VDD sky130_fd_sc_hd__inv_2
X_1912_ VSS VDD _1024_ core.ndc.rowon_out_n\[15\] _1331_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_8_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2892_ VSS VDD _0666_ _0785_ _0702_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1843_ VDD VSS _1324_ _1331_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_1774_ VDD VSS _1284_ _1095_ VSS VDD sky130_fd_sc_hd__buf_2
Xgenblk2\[11\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[11\] core.ndc.rowon_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2326_ VDD VSS _0349_ _0347_ _0348_ VSS VDD sky130_fd_sc_hd__and2_1
X_2257_ VSS VDD _0284_ _0286_ _0283_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_84_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2188_ VSS VDD core.cnb.next_average_sum_w\[1\] _0225_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_92_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1976__A1 _1208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[7\].buf_n_rown_A core.ndc.row_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_rowoff_n[0] core.pdc.rowoff_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_35 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_305 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_75_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_124_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1664__B1 _1035_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_393 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1719__A1 _1064_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1490_ VDD VSS core.cnb.data_register_r\[7\] _1050_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_3160_ VSS VDD net63 core.osr.next_result_w\[0\] net81 core.osr.result_r\[0\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_3091_ VSS VDD _0975_ _0976_ _0691_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2111_ VSS VDD _1413_ _0164_ _1101_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2042_ VSS VDD _0089_ _0123_ _1279_ VSS VDD sky130_fd_sc_hd__nand2_1
Xgenblk1\[28\].buf_n_coln VDD VSS core.ndc.col_out_n\[28\] nmatrix_col_core_n_buffered\[28\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_50_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xobstruction1 VDD VSS scboundary
X_2944_ VSS VDD _0834_ _0836_ _0835_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1958__A1 _1057_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2875_ VSS VDD _0685_ _0695_ _0769_ _0693_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1826_ VSS VDD core.cnb.data_register_r\[9\] _1071_ _1317_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1757_ VSS VDD _1272_ _1225_ _1273_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1688_ VSS VDD _1074_ _1224_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA_nmat_col[7] core.ndc.col_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2309_ VSS VDD _0326_ _0333_ _0332_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_85_422 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2438__A2 _1340_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1511__A _1037_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2610__A2 core.osr.next_result_w\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[30\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[30\] core.ndc.col_out_n\[30\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2061__B _1093_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_102 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_95_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_91_414 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_56_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2062__B1 _1075_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2252__A core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2660_ VSS VDD _0561_ _0041_ _0564_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1611_ VDD VSS _1159_ _1158_ VSS VDD sky130_fd_sc_hd__inv_2
X_2591_ VSS VDD _0030_ _0506_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1542_ VDD VSS _1098_ _1097_ VSS VDD sky130_fd_sc_hd__inv_2
X_1473_ VDD VSS _1032_ _1033_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_10_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3143_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0033_ net79 core.cnb.result_out\[11\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_3074_ VSS VDD _0960_ _0959_ _0958_ _0918_ _1312_ VSS VDD sky130_fd_sc_hd__a211o_1
X_2025_ VSS VDD _0101_ _0112_ _1093_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2927_ VSS VDD _0815_ _0726_ _0819_ _0818_ VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__1985__B _1275_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[8\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[8\] core.ndc.rowon_out_n\[8\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2858_ VSS VDD _0727_ _0752_ _0753_ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk2\[1\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[1\] core.pdc.row_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1809_ VSS VDD net14 _1301_ _1302_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2789_ VDD VSS _0685_ _0684_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1506__A _1034_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1619__A0 _1161_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1416__A core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2712_ VDD VSS _0348_ _0347_ _0528_ _0611_ VSS VDD sky130_fd_sc_hd__a21o_1
X_2643_ VSS VDD _0039_ _0548_ _0540_ _0547_ _0549_ VSS VDD sky130_fd_sc_hd__a31o_1
X_2574_ VSS VDD _0492_ _0494_ _0493_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1525_ VSS VDD _1083_ _1076_ _1078_ _1080_ _1082_ VSS VDD sky130_fd_sc_hd__o211a_1
X_1456_ VSS VDD _1019_ _1020_ _0983_ VSS VDD sky130_fd_sc_hd__nor2_2
X_3126_ VSS VDD clknet_2_2__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[4\]
+ net89 core.cnb.average_counter_r\[4\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_27_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_3057_ VSS VDD _0942_ _0944_ _0902_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2008_ VSS VDD _1131_ _0098_ _0099_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_50_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2026__B1 _1064_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1552__A2 _1096_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_76_46 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_132_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2017__A0 _1137_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2290_ VSS VDD core.osr.result_r\[9\] _0315_ core.cnb.result_out\[9\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_110_146 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2143__C core.cnb.sampled_avg_control_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2626_ VSS VDD core.osr.next_result_w\[8\] _0534_ _0533_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2440__A _1342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2557_ VSS VDD _0438_ _0480_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2488_ VDD VSS core.cnb.next_conv_finished_w _0434_ VSS VDD sky130_fd_sc_hd__inv_2
X_1508_ VDD VSS _1066_ _1065_ VSS VDD sky130_fd_sc_hd__inv_2
X_1439_ VDD VSS _1003_ _1002_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_87_347 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3109_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0009_ net90 core.cnb.shift_register_r\[7\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_15_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_59 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_483 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2334__B _0241_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1525__A2 _1078_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xinput13 VSS VDD net13 config_1_in[5] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1790_ VDD VSS _1294_ _1109_ VSS VDD sky130_fd_sc_hd__inv_2
Xinput24 VSS VDD config_2_in[15] net24 VSS VDD sky130_fd_sc_hd__clkbuf_2
Xinput35 VSS VDD net35 start_conversion_in VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2411_ VDD VSS _0418_ core.osr.next_sample_count_w\[6\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2342_ VSS VDD _0360_ _0363_ _0362_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_96_144 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2273_ VDD VSS _0300_ _0299_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1604__A _1092_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_269 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1988_ VSS VDD _0084_ _0085_ _1235_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2170__A _0210_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2609_ VSS VDD _1009_ _1018_ _0520_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA_nmat_col[29] core.ndc.col_out\[29\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1514__A net15 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1691__A1 _1224_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_98 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1424__A _0983_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1682__A1 _1078_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2960_ VSS VDD _0850_ _0852_ _0851_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1911_ VSS VDD _1378_ _1379_ _1369_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2891_ VSS VDD _0784_ _0783_ _0470_ VSS VDD sky130_fd_sc_hd__nand2_2
X_1842_ VSS VDD _1325_ _1328_ _1330_ core.pdc.row_out_n\[4\] VSS VDD sky130_fd_sc_hd__o21a_1
XANTENNA__3086__A _1342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1773_ VDD VSS core.ndc.col_out_n\[24\] core.ndc.col_out\[24\] VSS VDD sky130_fd_sc_hd__clkinv_2
Xgenblk2\[6\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[6\] core.pdc.row_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_69_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2325_ VSS VDD _0348_ core.cnb.result_out\[11\] _0255_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__3130__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2256_ VSS VDD _0285_ _0283_ _0284_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_27_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2187_ VSS VDD _0225_ _0224_ _0223_ _0209_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_53_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1988__B _1235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2165__A _0208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_43_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_68_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_124_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_sample sample_nmatrix_cgen VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1664__A1 _1075_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_129_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk1\[1\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[1\] core.pdc.col_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_3090_ VSS VDD _0972_ _0975_ _0974_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2110_ VSS VDD _1411_ _0163_ _1177_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_12_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2041_ VDD VSS core.pdc.col_out_n\[13\] core.pdc.col_out\[13\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2943_ VDD VSS _0835_ _0829_ VSS VDD sky130_fd_sc_hd__inv_2
Xobstruction2 VDD VSS scboundary
X_2874_ VSS VDD _0662_ _0664_ _0768_ _0767_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_88_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1825_ VDD VSS core.pdc.rowoff_out_n\[8\] _1316_ VSS VDD sky130_fd_sc_hd__buf_2
X_1756_ VSS VDD _1110_ _1272_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1687_ VDD VSS core.ndc.col_out_n\[11\] core.ndc.col_out\[11\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1591__B1 _1088_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col[6] core.ndc.col_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2308_ VDD VSS _0332_ _0330_ VSS VDD sky130_fd_sc_hd__inv_2
X_2239_ VDD VSS _0251_ core.cnb.result_out\[3\] _0269_ _0270_ VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_53_342 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_16 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2623__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[3\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[3\] core.ndc.row_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_134_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_119_75 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_79_35 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_102_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_79_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_114 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_input22_A config_2_in[13] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_404 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_91_426 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_56_180 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2062__A1 _1064_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1610_ VSS VDD _1158_ _1073_ _1119_ VSS VDD sky130_fd_sc_hd__or2_1
X_2590_ VSS VDD _0506_ core.cnb.result_out\[8\] _0480_ _0505_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1541_ VSS VDD _1047_ _1097_ _1057_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1472_ VSS VDD core.cnb.data_register_r\[8\] _1032_ net15 VSS VDD sky130_fd_sc_hd__nor2_2
X_3142_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0032_ net81 core.cnb.result_out\[10\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3073_ VDD VSS _0958_ _0831_ _0856_ _0959_ VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__2427__B core.pdc.rowoff_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2024_ VDD VSS _0083_ _1409_ _1208_ _0111_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_50_389 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2926_ VSS VDD _0649_ _0817_ _0818_ _0724_ VSS VDD sky130_fd_sc_hd__nand3_2
X_2857_ VSS VDD _0743_ _0745_ _0752_ _0751_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1808_ VDD VSS _1301_ core.cnb.data_register_r\[11\] VSS VDD sky130_fd_sc_hd__inv_2
X_2788_ VSS VDD _0680_ _0683_ _0684_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1739_ VDD VSS core.ndc.col_out\[18\] core.ndc.col_out_n\[18\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_49_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1522__A _1079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_65_59 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_121_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2044__A1 _1161_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2072__B _1275_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1555__B1 _1088_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_106 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2711_ VSS VDD _0607_ _0610_ _0609_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2642_ VDD VSS _0393_ _0542_ core.osr.next_result_w\[1\] _0549_ net49 VSS VDD sky130_fd_sc_hd__a22o_1
X_2573_ VSS VDD _0489_ _0493_ _1200_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1607__A _1101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1524_ VDD VSS _1081_ _1082_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_1455_ VDD VSS _1019_ _1018_ VSS VDD sky130_fd_sc_hd__inv_2
X_3125_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[3\]
+ net89 core.cnb.average_counter_r\[3\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3056_ VSS VDD _0689_ _0943_ _0058_ _1312_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_35_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2007_ VSS VDD _1389_ _1229_ _1161_ _0098_ VSS VDD sky130_fd_sc_hd__mux2_2
XANTENNA__2026__A1 _1224_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_186 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2909_ VSS VDD _0798_ _0801_ _0800_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1517__A _1074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1537__B1 _1075_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_111 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout72_A net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_404 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_26_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_92_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2017__A1 _1133_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_110_114 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[10\].buf_p_rown_A core.pdc.row_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2625_ VSS VDD _1000_ _0533_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2556_ VSS VDD _0477_ _0479_ _0478_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2487_ VSS VDD _0220_ _0434_ core.cnb.is_holding_result_w VSS VDD sky130_fd_sc_hd__nand2_1
X_1507_ VSS VDD core.cnb.data_register_r\[4\] _1065_ _1044_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1438_ VSS VDD _1000_ _1002_ _0989_ VSS VDD sky130_fd_sc_hd__nor2_2
XANTENNA__2168__A _0210_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3108_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0008_ net90 core.cnb.shift_register_r\[6\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3039_ VSS VDD _0856_ _0927_ _0924_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_51_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_102_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_127_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_87_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk1\[6\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[6\] core.pdc.col_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2078__A _0065_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1710__A _1117_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput14 VDD VSS net14 config_1_in[6] VSS VDD sky130_fd_sc_hd__buf_2
Xinput25 VSS VDD net25 config_2_in[1] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2410_ VSS VDD _1021_ _0417_ _0416_ _0418_ VSS VDD sky130_fd_sc_hd__or3b_1
X_2341_ VSS VDD _0355_ _0362_ _0361_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2272_ _0299_ _0297_ _0298_ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA__3091__B _0691_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3183__RESET_B net86 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1987_ VSS VDD _0084_ _1036_ _1053_ _1390_ _0083_ VSS VDD sky130_fd_sc_hd__a31o_1
Xgenblk2\[8\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[8\] core.ndc.row_out_n\[8\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2608_ VSS VDD _0518_ _0519_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2539_ VSS VDD _0188_ _0463_ _0235_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col[28] core.ndc.col_out\[28\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2626__A core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_384 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_113_77 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_138_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_98_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1705__A core.ndc.col_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2536__A _0438_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1682__A2 _1135_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1910_ VSS VDD _1355_ _1378_ _1342_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_63_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2890_ VSS VDD _0759_ _0783_ _0770_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1841_ VSS VDD _1329_ _1330_ _1302_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2271__A core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3086__B _0799_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1772_ VSS VDD core.ndc.col_out_n\[24\] _1283_ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xgenblk1\[3\].buf_n_coln VDD VSS core.ndc.col_out_n\[3\] nmatrix_col_core_n_buffered\[3\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_2324_ VSS VDD _0345_ _0271_ _0347_ _0346_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_69_134 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2255_ VSS VDD _0277_ _0284_ _0273_ VSS VDD sky130_fd_sc_hd__nand2_1
Xpmat_sample_buf_n VSS VDD pmat_sample_switch_n_buffered core.cnb.enable_loop_out
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2186_ VDD VSS core.cnb.average_sum_r\[0\] core.cnb.comparator_in core.cnb.average_sum_r\[1\]
+ _0224_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__2622__A1 _0254_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_119 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_88_410 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_108_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_88_454 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__3162__D core.osr.next_result_w\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_351 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_74 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2613__B2 core.osr.next_result_w\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_33_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2129__B1 _1121_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2040_ VSS VDD core.pdc.col_out_n\[13\] _0122_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_47_373 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2942_ VSS VDD _0753_ _0832_ _0834_ _0833_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2873_ VDD VSS _0767_ _0708_ _0766_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_90_90 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1824_ VDD VSS _1316_ _1302_ VSS VDD sky130_fd_sc_hd__inv_2
X_1755_ VDD VSS core.ndc.col_out\[21\] core.ndc.col_out_n\[21\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1591__A1 _1105_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1686_ VSS VDD _1223_ core.ndc.col_out_n\[11\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA_nmat_col[5] core.ndc.col_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2307_ VSS VDD _0326_ _0331_ _0330_ VSS VDD sky130_fd_sc_hd__or2b_1
X_2238_ VSS VDD _0269_ _0268_ _0267_ _0988_ VSS VDD sky130_fd_sc_hd__and3_1
X_2169_ VSS VDD core.cnb.next_average_counter_w\[1\] _0211_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_72_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_110_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_119_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_119_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_134_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_79_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1582__A1 _1079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_95_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_input15_A config_1_in[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1702__B _1235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_61 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2598__B1 _1022_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3120__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3011__A1 _1053_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1540_ VDD VSS _1096_ _1095_ VSS VDD sky130_fd_sc_hd__buf_2
X_1471_ VSS VDD core.ndc.rowoff_out_n\[0\] core.ndc.row_out_n\[0\] core.ndc.rowon_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_3141_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0031_ net77 core.cnb.result_out\[9\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_54_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col_n[29] nmatrix_col_core_n_buffered\[29\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3072_ VSS VDD _0958_ _0833_ _0726_ _0910_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_54_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2023_ VDD VSS _0110_ _0108_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_50_302 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2925_ VSS VDD _0659_ _0816_ _0699_ _0817_ VSS VDD sky130_fd_sc_hd__nor3_1
X_2856_ VDD VSS _0751_ _0750_ VSS VDD sky130_fd_sc_hd__inv_2
X_1807_ VSS VDD core.cnb.data_register_r\[8\] _1300_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2787_ VSS VDD _0640_ _0683_ _0682_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1738_ VSS VDD _1035_ _1231_ _1260_ _1259_ core.ndc.col_out_n\[18\] _1261_ VSS VDD
+ sky130_fd_sc_hd__o221a_2
X_1669_ VSS VDD _1209_ _1197_ _1054_ _1208_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A config_1_in[14] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1803__A core.ndc.col_out\[31\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1867__A2 _1325_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2634__A _0983_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3143__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_30_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1555__A1 _1037_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_30_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_122_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1432__B _0995_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2710_ VDD VSS _0609_ _0608_ VSS VDD sky130_fd_sc_hd__inv_2
X_2641_ VSS VDD _0548_ _0537_ core.osr.next_result_w\[3\] VSS VDD sky130_fd_sc_hd__or2_1
X_2572_ VSS VDD _0492_ _1200_ _0489_ VSS VDD sky130_fd_sc_hd__or2_1
X_1523_ VSS VDD core.cnb.data_register_r\[7\] _1081_ _1058_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1454_ VSS VDD _1018_ _1006_ _1017_ VSS VDD sky130_fd_sc_hd__nand2_2
XANTENNA__1623__A _1128_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_sample_buf_A net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3124_ VSS VDD clknet_2_2__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[2\]
+ net89 core.cnb.average_counter_r\[2\] VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3055_ VSS VDD _0905_ _0943_ _0942_ _0781_ _0936_ VSS VDD sky130_fd_sc_hd__o211ai_1
X_2006_ VDD VSS core.pdc.col_out_n\[8\] core.pdc.col_out\[8\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_50_110 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2908_ VSS VDD _0799_ _0800_ _0796_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2982__B1 _1114_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2839_ VSS VDD _0733_ _0730_ _0734_ _0731_ VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__1537__A1 _1064_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_123 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_116_55 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout65_A net66 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk2\[4\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[4\] core.ndc.rowon_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_92_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_rowon_n[1] nmatrix_rowon_core_n_buffered\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[8\].buf_n_coln VDD VSS core.ndc.col_out_n\[8\] nmatrix_col_core_n_buffered\[8\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_110_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_110_126 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3189__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2624_ VSS VDD _0037_ _0531_ _0529_ _0532_ VSS VDD sky130_fd_sc_hd__a21bo_1
XANTENNA__1618__A _1163_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2555_ VSS VDD _0474_ _0478_ core.cnb.pswitch_out\[1\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2486_ VDD VSS _0001_ sample_nmatrix_cgen VSS VDD sky130_fd_sc_hd__inv_2
X_1506_ VDD VSS _1064_ _1034_ VSS VDD sky130_fd_sc_hd__buf_2
X_1437_ VSS VDD _1000_ _1001_ core.osr.osr_mode_r\[0\] VSS VDD sky130_fd_sc_hd__nor2_2
X_3107_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0007_ net88 core.cnb.shift_register_r\[5\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_55_235 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3038_ VSS VDD _0925_ _0926_ _0475_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2184__A core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1758__A1 _1121_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1758__B2 _1125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1528__A _1079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_87_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1710__B _1060_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput15 VDD VSS net15 config_1_in[7] VSS VDD sky130_fd_sc_hd__buf_2
Xinput26 VSS VDD net26 config_2_in[2] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2340_ VDD VSS _0361_ core.osr.result_r\[13\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_96_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2271_ VSS VDD core.cnb.result_out\[7\] _0298_ core.osr.result_r\[7\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_78_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1986_ VDD VSS _0083_ _1206_ VSS VDD sky130_fd_sc_hd__inv_2
X_2607_ VDD VSS _0518_ _1001_ VSS VDD sky130_fd_sc_hd__inv_2
X_2538_ VSS VDD _0178_ _0222_ _0462_ _0187_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_87_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2469_ VDD VSS core.ndc.rowoff_out_n\[15\] _0432_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_69_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_113_23 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_113_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1530__B _1085_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_22_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1840_ VSS VDD _1326_ _1023_ _1329_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_8_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1771_ VSS VDD _1283_ _1282_ _1281_ _1280_ VSS VDD sky130_fd_sc_hd__and3_1
X_2323_ VSS VDD _0338_ _0328_ _0346_ _0343_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2254_ VDD VSS _0283_ _0281_ _0282_ VSS VDD sky130_fd_sc_hd__and2_1
X_2185_ VSS VDD _0218_ core.cnb.average_sum_r\[1\] _0222_ _0223_ VSS VDD sky130_fd_sc_hd__or3b_1
XANTENNA__1631__A _1072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1969_ VDD VSS _0070_ _0069_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1806__A core.pdc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_88_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_477 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1649__B1 _1082_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1541__A _1047_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_56_385 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2091__B _1101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2129__A1 _1126_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_385 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_74_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2941_ VDD VSS _0833_ _0806_ VSS VDD sky130_fd_sc_hd__inv_2
X_2872_ VSS VDD _0765_ _0766_ _0635_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1823_ VSS VDD _1315_ core.pdc.row_out_n\[1\] _1307_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1754_ VSS VDD _1271_ core.ndc.col_out_n\[21\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1591__A2 _1104_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1685_ VSS VDD _1223_ _1222_ _1219_ _1218_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA_nmat_col[4] core.ndc.col_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2306_ VSS VDD _0327_ _0329_ _0330_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2237_ VSS VDD _0268_ _0266_ _0263_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__2457__A core.ndc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2168_ VSS VDD _0211_ _0191_ _0182_ _0210_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_53_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2099_ VDD VSS _0081_ _1173_ core.pdc.col_out\[25\] _0079_ _1096_ _0157_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1536__A _1091_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1582__A2 _1113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_63_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_491 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2598__A1 _1328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[12\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[12\] core.pdc.rowon_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_125_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_60_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1470_ VSS VDD _1031_ core.ndc.rowon_out_n\[0\] _1030_ VSS VDD sky130_fd_sc_hd__nand2_4
X_3140_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0030_ net81 core.cnb.result_out\[8\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA_nmat_col_n[28] nmatrix_col_core_n_buffered\[28\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3071_ VSS VDD _0936_ _0957_ _0956_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2022_ VDD VSS core.pdc.col_out_n\[10\] core.pdc.col_out\[10\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_62_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_genblk2\[8\].buf_p_rown_A core.pdc.row_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2924_ VDD VSS _0816_ _0645_ VSS VDD sky130_fd_sc_hd__inv_2
X_2855_ VSS VDD _0454_ _0749_ _0750_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1806_ VSS VDD core.pdc.rowon_out_n\[0\] core.pdc.row_out_n\[0\] core.pdc.rowoff_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2786_ VSS VDD _0681_ _0659_ _0682_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA_genblk2\[13\].buf_p_rowonn_A core.pdc.rowon_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1737_ VSS VDD _1261_ _1074_ _1204_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_131_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1668_ VSS VDD _1206_ _1207_ _1208_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1599_ VDD VSS _1149_ _1148_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_105_35 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3168__D core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_225 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2640_ VSS VDD _0544_ _0545_ _0547_ _0546_ VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__2560__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2571_ VSS VDD _0025_ _0439_ _0489_ _0490_ _0491_ VSS VDD sky130_fd_sc_hd__o31a_1
X_1522_ VDD VSS _1080_ _1079_ VSS VDD sky130_fd_sc_hd__inv_2
X_1453_ VDD VSS _1017_ _1016_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_87_509 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_113_124 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3123_ VSS VDD clknet_2_2__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[1\]
+ net88 core.cnb.average_counter_r\[1\] VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_27_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3054_ VSS VDD _0941_ _0942_ _0905_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2005_ VSS VDD _1035_ _0072_ _0094_ _1126_ core.pdc.col_out_n\[8\] _0097_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2907_ VDD VSS _0784_ _0799_ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__2470__A core.pdc.row_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2838_ VSS VDD _0638_ _0658_ _0733_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2769_ VSS VDD _0662_ _0664_ _0665_ _0658_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__2734__A1 core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_116_67 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3110__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_66 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout58_A net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_26_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_92_37 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_494 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_rowon_n[0] nmatrix_rowon_core_n_buffered\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_266 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_501 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[9\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[9\] core.pdc.rowon_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_32_111 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_82_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2623_ VSS VDD _0394_ _0532_ net47 VSS VDD sky130_fd_sc_hd__nand2_1
X_2554_ VSS VDD _0477_ core.cnb.pswitch_out\[1\] _0474_ VSS VDD sky130_fd_sc_hd__or2_1
X_1505_ VDD VSS core.ndc.col_out\[0\] core.ndc.col_out_n\[0\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_99_133 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1634__A _1179_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2485_ VSS VDD sample_pmatrix_cgen _0000_ VSS VDD sky130_fd_sc_hd__inv_1
X_1436_ VDD VSS _1000_ _0994_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__3133__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_101_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3106_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0006_ net88 core.cnb.shift_register_r\[4\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_83_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3037_ VSS VDD _0831_ _0925_ _0924_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_62_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1809__A net14 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1758__A2 _1193_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1528__B _1085_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_88 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_309 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_36_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xinput16 VSS VDD net16 config_1_in[8] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput27 VSS VDD net27 config_2_in[3] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA_genblk1\[1\].buf_n_coln_A core.ndc.col_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_7 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_6 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2270_ VSS VDD core.cnb.result_out\[7\] core.osr.result_r\[7\] _0297_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_20_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1985_ VSS VDD _0081_ _0082_ _1275_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2606_ VSS VDD _1003_ _0517_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__3121__RESET_B net86 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2537_ VSS VDD _0460_ _0461_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2468_ VDD VSS _0432_ core.ndc.row_out_n\[15\] core.ndc.rowon_out_n\[15\] VSS VDD
+ sky130_fd_sc_hd__and2_1
XFILLER_87_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1419_ VDD VSS _0982_ _0983_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_2399_ VSS VDD core.osr.sample_count_r\[4\] _0405_ _0409_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_56_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_113_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1539__A _1072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3179__CLK net58 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_22_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2864__B1 core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1770_ VSS VDD _1172_ _1282_ _1095_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2322_ VSS VDD _0339_ _0345_ _0344_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2253_ VSS VDD core.cnb.result_out\[5\] _0282_ core.osr.result_r\[5\] VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_sample_n_in net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2184_ VDD VSS _0222_ core.cnb.comparator_in VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2727__B _1002_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_515 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2462__B core.ndc.rowon_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1968_ VSS VDD _0069_ _1105_ _1104_ _1403_ _1088_ VSS VDD sky130_fd_sc_hd__a31o_1
X_1899_ VDD VSS core.pdc.rowon_out_n\[3\] _1371_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1806__B core.pdc.rowoff_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_75_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1649__A1 _1128_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1541__B _1057_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_397 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2940_ VSS VDD _0809_ _0819_ _0832_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2871_ VSS VDD core.cnb.shift_register_r\[4\] _0705_ _0765_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1822_ VSS VDD _1311_ _1314_ _1315_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_90_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_128_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1753_ VSS VDD _1271_ _1209_ _1034_ _1139_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1684_ VSS VDD _1221_ _1222_ _1177_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col[3] core.ndc.col_out\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2305_ VDD VSS _0329_ _0328_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1642__A _1117_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2236_ VSS VDD _0263_ _0267_ _0266_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2457__B core.ndc.rowon_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2167_ VSS VDD _0210_ core.cnb.next_average_counter_w\[0\] core.cnb.average_counter_r\[0\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2098_ VSS VDD _0065_ _0115_ _0157_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2473__A core.pdc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1567__B1 _1075_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_134_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1536__B _1093_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_71_120 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_125_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3070_ VSS VDD _0904_ _0948_ _0956_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2021_ VSS VDD _1064_ _0076_ _0106_ _1224_ core.pdc.col_out_n\[10\] _0109_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XFILLER_47_194 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2923_ VSS VDD _0750_ _0814_ _0815_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2854_ VSS VDD _0748_ _0749_ _0649_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1805_ VSS VDD _1030_ core.pdc.rowoff_out_n\[0\] _1027_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2785_ VSS VDD _0644_ _0681_ _0642_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_116_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1736_ VDD VSS _1260_ _1124_ VSS VDD sky130_fd_sc_hd__inv_2
X_1667_ VSS VDD _1113_ _1057_ _1207_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_131_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1598_ VSS VDD _1148_ _1147_ _1077_ _1146_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_105_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2219_ VSS VDD _0251_ _0252_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__2277__A1 core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3199_ VSS VDD net64 core.osr.next_sample_count_w\[7\] net77 core.osr.sample_count_r\[7\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_121_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_121_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_81_39 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1547__A _1078_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_input20_A config_2_in[11] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_237 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2570_ VSS VDD _0491_ core.cnb.result_out\[3\] _0461_ VSS VDD sky130_fd_sc_hd__or2_1
X_1521_ VSS VDD _1079_ _1044_ _1055_ VSS VDD sky130_fd_sc_hd__nand2_2
X_1452_ VDD VSS _1003_ _1007_ _1016_ _1010_ _1012_ _1015_ VSS VDD sky130_fd_sc_hd__a221o_1
XFILLER_113_136 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3122_ VDD VSS core.cnb.average_counter_r\[0\] net88 core.cnb.next_average_counter_w\[0\]
+ clknet_2_2__leaf_clk_dig_dummy VSS VDD sky130_fd_sc_hd__dfstp_1
X_3053_ VSS VDD _0937_ _0941_ _0940_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2004_ VSS VDD _0096_ _0097_ _1284_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2431__B2 core.ndc.row_bottotop_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2906_ VSS VDD _0795_ _0798_ _0797_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2470__B core.pdc.rowon_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2837_ VSS VDD _0729_ _0730_ _0732_ _0731_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2768_ VSS VDD _0640_ _0647_ _0664_ _0663_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2699_ VSS VDD _0596_ _0597_ _0599_ _0598_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1719_ VSS VDD _1075_ _1246_ _1183_ _1064_ core.ndc.col_out_n\[15\] _1248_ VSS VDD
+ sky130_fd_sc_hd__o221a_2
XANTENNA__1942__A0 _1067_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_132_34 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_cgen_start_conv_in net35 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_92_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1724__B _1213_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk1\[10\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[10\] core.pdc.col_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_2_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_513 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2555__B core.cnb.pswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2622_ VDD VSS _0530_ _0254_ _1018_ _0531_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_2553_ VSS VDD _0476_ _0461_ core.cnb.result_out\[0\] _0474_ _0022_ VSS VDD sky130_fd_sc_hd__o22a_1
X_1504_ VSS VDD core.ndc.col_out_n\[0\] _1063_ _1049_ _1035_ VSS VDD sky130_fd_sc_hd__o21a_2
X_2484_ VDD VSS core.cnb.enable_loop_out net55 VSS VDD sky130_fd_sc_hd__inv_2
X_1435_ VDD VSS _0999_ core.osr.sample_count_r\[4\] VSS VDD sky130_fd_sc_hd__inv_2
X_3105_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0005_ net88 core.cnb.shift_register_r\[3\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3036_ VDD VSS _0924_ _0923_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1650__A _1077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2465__B _1325_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_102_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_102_59 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2481__A core.pdc.row_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A net83 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk1\[16\].buf_n_coln_A core.ndc.col_out_n\[16\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput17 VSS VDD net17 config_1_in[9] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput28 VDD VSS net28 config_2_in[4] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xgenblk2\[0\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[0\] core.ndc.rowon_out_n\[0\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
Xgenblk2\[14\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[14\] core.pdc.row_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2566__A core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1984_ VSS VDD _0081_ _1112_ _1409_ _1118_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2605_ VDD VSS _0395_ _0516_ _0995_ _0034_ net38 VSS VDD sky130_fd_sc_hd__a22o_1
XANTENNA_nmat_col[25] core.ndc.col_out\[25\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1645__A _1187_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2536_ VDD VSS _0460_ _0438_ VSS VDD sky130_fd_sc_hd__inv_2
X_2467_ VSS VDD core.ndc.row_out_n\[14\] core.ndc.rowoff_out_n\[14\] core.ndc.rowon_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_genblk1\[6\].buf_p_coln_A core.pdc.col_out_n\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1418_ VDD VSS net11 net13 net12 _0982_ VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_87_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2398_ VDD VSS core.osr.next_sample_count_w\[3\] _0408_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_83_365 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3019_ VSS VDD _0804_ _0870_ _0907_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_51_251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2864__B2 _0758_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2833__B _0637_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__3123__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2321_ VDD VSS _0344_ _0343_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2552__B1 core.cnb.pswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2252_ VSS VDD _0281_ core.cnb.result_out\[5\] core.osr.result_r\[5\] VSS VDD sky130_fd_sc_hd__or2_1
X_2183_ VDD VSS core.cnb.comparator_in core.cnb.next_average_sum_w\[0\] _0221_ VSS
+ VDD sky130_fd_sc_hd__xor2_1
XFILLER_138_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1967_ VDD VSS _0068_ _1407_ VSS VDD sky130_fd_sc_hd__inv_2
X_1898_ VSS VDD _1370_ _1309_ _1371_ _1305_ VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_108_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_108_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk2\[11\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[11\] core.ndc.row_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_68_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2519_ VSS VDD _0451_ core.cnb.shift_register_r\[13\] _0219_ core.cnb.shift_register_r\[12\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_56_321 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_56_365 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_87 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2534__A0 core.cnb.sampled_avg_control_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_58_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2870_ VSS VDD _0702_ _0764_ _0763_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_71_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1821_ VDD VSS _1314_ _1313_ VSS VDD sky130_fd_sc_hd__inv_2
X_1752_ VDD VSS core.ndc.col_out_n\[20\] core.ndc.col_out\[20\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_1683_ VDD VSS _1221_ _1220_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col[2] core.ndc.col_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2304_ VSS VDD core.osr.result_r\[10\] _0328_ core.cnb.result_out\[10\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2235_ VDD VSS _0266_ _0264_ _0265_ VSS VDD sky130_fd_sc_hd__and2_1
X_2166_ VSS VDD _0209_ _0210_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__3169__CLK net66 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2097_ VDD VSS core.pdc.col_out_n\[24\] core.pdc.col_out\[24\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_62_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2999_ VSS VDD _0763_ _0888_ _0695_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1567__A1 _1064_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_298 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[15\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[15\] core.pdc.col_out_n\[15\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_71_132 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_69_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1743__A _1227_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2020_ VSS VDD _0108_ _0109_ _1093_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_90_441 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_463 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2922_ VSS VDD _0737_ _0811_ _0814_ _0813_ VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__1918__A _1381_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2853_ VSS VDD _0646_ _0673_ _0747_ _0748_ VSS VDD sky130_fd_sc_hd__nor3_1
X_1804_ VSS VDD core.pdc.rowon_out_n\[0\] _1025_ _1031_ VSS VDD sky130_fd_sc_hd__nand2_2
X_2784_ VDD VSS _0680_ _0679_ VSS VDD sky130_fd_sc_hd__inv_2
X_1735_ VSS VDD _1110_ _1259_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1637__B _1096_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1666_ VSS VDD _1206_ _1059_ _1052_ VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_131_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1597_ VSS VDD _1123_ _1147_ _1068_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2218_ VDD VSS _0251_ _0988_ VSS VDD sky130_fd_sc_hd__inv_2
X_3198_ VSS VDD net64 core.osr.next_sample_count_w\[6\] net77 core.osr.sample_count_r\[6\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2149_ VSS VDD _0193_ _0190_ _0192_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_53_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2484__A net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_30_99 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2268__A2 _0255_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_205 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_input13_A config_1_in[5] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_249 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1520_ VDD VSS _1078_ _1077_ VSS VDD sky130_fd_sc_hd__buf_2
X_1451_ VDD VSS core.osr.sample_count_r\[8\] _0992_ _1014_ _1015_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__2569__A _1395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1473__A _1032_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[12\].buf_n_coln VDD VSS core.ndc.col_out_n\[12\] nmatrix_col_core_n_buffered\[12\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_3121_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0021_ net86 core.cnb.sampled_avg_control_r\[2\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA__2259__A2 _0240_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_460 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3052_ VDD VSS _0940_ _0939_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_48_482 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2003_ VDD VSS _0096_ _0095_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__3186__RESET_B net85 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2905_ VDD VSS _0797_ _0796_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1648__A core.ndc.col_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2836_ VDD VSS _0731_ _0724_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_2767_ VSS VDD core.cnb.shift_register_r\[9\] _0633_ _0663_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2698_ VSS VDD core.osr.next_result_w\[14\] _0598_ _0535_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1718_ VSS VDD _1247_ _1248_ _1093_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_104_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2479__A core.pdc.rowon_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_rowon_n[12] nmatrix_rowon_core_n_buffered\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1649_ VDD VSS core.cnb.data_register_r\[7\] _1128_ _1082_ _1191_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA_genblk2\[4\].buf_p_rown_A core.pdc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input5_A config_1_in[12] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_132_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_41_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2186__A1 core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_393 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1740__B _1152_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_61 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2621_ VSS VDD _1009_ _0530_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2552_ VDD VSS _0475_ _0461_ core.cnb.pswitch_out\[0\] _0476_ VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__1915__B core.ndc.rowon_bottotop_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1503_ VDD VSS _1063_ _1062_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_99_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2483_ VDD VSS _0433_ core.pdc.rowoff_out_n\[15\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_1434_ VSS VDD _0996_ _0998_ core.osr.sample_count_r\[0\] VSS VDD sky130_fd_sc_hd__nand2_1
X_3104_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0004_ net88 core.cnb.shift_register_r\[2\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_83_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3035_ VSS VDD _0853_ _0923_ _0827_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_23_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_135 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2481__B core.pdc.rowon_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_499 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1612__B1 _1155_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2819_ VSS VDD _0692_ _0714_ _0713_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_11_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_127_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_127_79 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_39 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_330 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_36_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout63_A net66 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput18 VSS VDD net18 config_2_in[0] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput29 VDD VSS net29 config_2_in[5] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2566__B core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_322 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1983_ VSS VDD _0079_ _0080_ _1279_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2604_ VSS VDD _0279_ _1018_ _0516_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1645__B _1188_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2535_ VSS VDD _0021_ _0459_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2466_ VSS VDD core.ndc.row_out_n\[13\] core.ndc.rowoff_out_n\[13\] core.ndc.rowon_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
Xgenblk2\[5\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[5\] core.pdc.rowon_bottotop_n\[5\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_87_149 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1417_ VDD VSS core.cnb.pswitch_out\[0\] core.cnb.data_register_r\[0\] VSS VDD sky130_fd_sc_hd__inv_2
X_2397_ VDD VSS _0404_ _0403_ _0407_ _0408_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__2476__B core.pdc.rowon_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3018_ VSS VDD _0895_ _0879_ _0906_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_11_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_78_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_86_171 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2616__A2 _0395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1746__A core.ndc.col_out_n\[19\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[22\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[22\] core.pdc.col_out_n\[22\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2001__B1 _1053_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2320_ VSS VDD _0340_ _0342_ _0343_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2251_ VDD VSS _0280_ core.cnb.result_out\[5\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1481__A core.ndc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2182_ VSS VDD _0218_ _0220_ _0221_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_92_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1966_ VDD VSS core.pdc.col_out\[3\] core.pdc.col_out_n\[3\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_1897_ VSS VDD _1338_ _1370_ _1369_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_108_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2518_ VSS VDD _0013_ _0450_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_88_425 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2487__A _0220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2449_ VDD VSS core.pdc.rowoff_out_n\[5\] _1369_ _1384_ core.ndc.rowon_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_84_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_56_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_56_377 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_99 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2534__A1 net10 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_58_52 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_0__leaf_clk_dig_dummy
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xgenblk1\[17\].buf_n_coln VDD VSS core.ndc.col_out_n\[17\] nmatrix_col_core_n_buffered\[17\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_47_300 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_355 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_74_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1820_ VSS VDD _1313_ core.cnb.data_register_r\[9\] _1022_ _1312_ VSS VDD sky130_fd_sc_hd__and3_1
X_1751_ VSS VDD core.ndc.col_out_n\[20\] _1270_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1682_ VSS VDD _1135_ _1078_ _1220_ _1137_ VSS VDD sky130_fd_sc_hd__a21oi_2
XANTENNA_nmat_col[1] core.ndc.col_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2303_ VSS VDD core.osr.result_r\[10\] core.cnb.result_out\[10\] _0327_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1923__B core.ndc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2234_ VSS VDD core.cnb.result_out\[3\] _0265_ core.osr.result_r\[3\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2165_ VDD VSS _0209_ _0208_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_93_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2096_ VDD VSS _0092_ _1275_ core.pdc.col_out\[24\] _0087_ _1102_ _0156_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2998_ VSS VDD _0884_ _0887_ _0877_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1949_ VDD VSS _1403_ _1389_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_135_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3113__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_288 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_56_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_450 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_71_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_100_71 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_60_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_125_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col_n[25] nmatrix_col_core_n_buffered\[25\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_85_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2921_ VSS VDD _0812_ _0730_ _0813_ _0724_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2852_ VSS VDD _0633_ _0747_ _0746_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1803_ VDD VSS core.ndc.col_out_n\[31\] core.ndc.col_out\[31\] VSS VDD sky130_fd_sc_hd__inv_2
X_2783_ VSS VDD core.cnb.shift_register_r\[15\] _0678_ _0679_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1734_ VDD VSS core.ndc.col_out\[17\] core.ndc.col_out_n\[17\] VSS VDD sky130_fd_sc_hd__inv_2
X_1665_ VDD VSS core.ndc.col_out\[9\] core.ndc.col_out_n\[9\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__3136__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1596_ VDD VSS _1146_ _1145_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_131_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1653__B _1104_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2217_ VSS VDD _0239_ _0248_ _0250_ _0243_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_38_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3197_ VSS VDD net64 core.osr.next_sample_count_w\[5\] net80 core.osr.sample_count_r\[5\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2148_ VSS VDD _0192_ _0184_ _0191_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_121_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2079_ VDD VSS _1102_ _0108_ core.pdc.col_out\[20\] _1125_ _0146_ _0147_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2434__B1 _1328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout93_A net94 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_217 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1450_ VSS VDD _0986_ _1014_ _1013_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3120_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0020_ net85 core.cnb.sampled_avg_control_r\[1\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3051_ VSS VDD _0938_ _0939_ _0893_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_48_494 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2002_ VSS VDD _1082_ _1403_ _1191_ _0095_ VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_50_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2904_ VSS VDD _0648_ _0796_ _0763_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2835_ VSS VDD _0660_ _0730_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2766_ VSS VDD _0660_ _0662_ _0661_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2697_ VSS VDD core.osr.next_result_w\[16\] _0597_ _0533_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1717_ VDD VSS _1247_ _1070_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2479__B core.pdc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1648_ VDD VSS core.ndc.col_out\[8\] core.ndc.col_out_n\[8\] VSS VDD sky130_fd_sc_hd__inv_2
X_1579_ VDD VSS _1130_ _1125_ _1106_ _1121_ _1124_ core.ndc.col_out\[4\] VSS VDD sky130_fd_sc_hd__a221o_2
XANTENNA__2495__A _0208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xgenblk1\[27\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[27\] core.pdc.col_out_n\[27\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_89_361 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_66_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_66_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_82_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2620_ VSS VDD _0527_ _0529_ _0528_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2551_ VSS VDD _0472_ _0475_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_2482_ VDD VSS _0433_ core.pdc.row_out_n\[15\] core.pdc.rowon_out_n\[15\] VSS VDD
+ sky130_fd_sc_hd__and2_1
X_1502_ VSS VDD _1053_ _1061_ _1062_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1433_ VSS VDD _0997_ core.osr.sample_count_r\[0\] _0996_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_101_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3103_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0003_ net85 core.cnb.is_holding_result_w
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_3034_ VSS VDD _0915_ _0921_ _0922_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_23_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1612__A1 _1152_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2818_ VSS VDD _0697_ _0704_ _0713_ _0712_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2749_ VSS VDD core.cnb.shift_register_r\[14\] _0645_ core.cnb.shift_register_r\[15\]
+ VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_11_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_127_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_100_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_342 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1569__A _1101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput19 VDD VSS net19 config_2_in[10] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2566__C _1076_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_345 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_378 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1842__A1 _1325_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1479__A net15 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1982_ VDD VSS _0079_ _0066_ VSS VDD sky130_fd_sc_hd__inv_2
Xgenblk1\[24\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[24\] core.ndc.col_out_n\[24\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2603_ VSS VDD _0033_ _0515_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2534_ VSS VDD _0459_ net10 net54 core.cnb.sampled_avg_control_r\[2\] VSS VDD sky130_fd_sc_hd__mux2_1
X_2465_ VSS VDD _1338_ core.ndc.rowoff_out_n\[12\] _1325_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2396_ VSS VDD _0394_ _0407_ _0406_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1416_ VDD VSS core.cnb.pswitch_out\[1\] core.cnb.data_register_r\[1\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1661__B _1202_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3017_ VDD VSS _0905_ _0904_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2086__A1 _0101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2086__B2 _1096_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1833__A1 core.pdc.rowoff_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3170__RESET_B net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_286 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_63_20 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3026__B1 _1117_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[0\].buf_n_rowonn_A core.ndc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1588__A0 _1133_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_132 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_genblk1\[12\].buf_n_coln_A core.ndc.col_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2250_ VDD VSS core.osr.next_result_w\[4\] _0279_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1762__A _1187_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_26_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1481__B _1040_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2577__B _1114_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2181_ VDD VSS _0220_ _0219_ VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1512__A0 _1067_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1965_ VDD VSS _1121_ _1411_ core.pdc.col_out\[3\] _1125_ _1413_ _0067_ VSS VDD sky130_fd_sc_hd__a221o_1
XANTENNA__1579__B1 _1106_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2532__S net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1896_ VDD VSS _1369_ _1362_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_2517_ VSS VDD _0450_ core.cnb.shift_register_r\[12\] _0444_ core.cnb.shift_register_r\[11\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_2448_ VSS VDD _1336_ _1385_ core.ndc.rowon_out_n\[9\] core.pdc.rowon_bottotop_n\[5\]
+ VSS VDD sky130_fd_sc_hd__a21oi_2
X_2379_ VSS VDD _1020_ _0393_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_83_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2008__A _1131_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_58_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_312 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_114_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_74_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_130_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1757__A _1272_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1750_ VSS VDD _1270_ _1269_ _1268_ _1267_ VSS VDD sky130_fd_sc_hd__and3_1
X_1681_ VSS VDD _1212_ _1219_ _1173_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col[0] core.ndc.col_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_analog_in ANTENNA_nmat_analog_in/DIODE VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2302_ VSS VDD _0323_ _0326_ _0325_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2233_ VSS VDD _0264_ core.cnb.result_out\[3\] core.osr.result_r\[3\] VSS VDD sky130_fd_sc_hd__or2_1
X_2164_ VSS VDD _0207_ _0208_ _0204_ VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_93_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2095_ VSS VDD _0065_ _0135_ _0156_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1667__A _1113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2997_ VSS VDD _0056_ _0885_ _0781_ _0884_ _0886_ VSS VDD sky130_fd_sc_hd__a31o_1
X_1948_ VDD VSS core.pdc.col_out_n\[1\] core.pdc.col_out\[1\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_1879_ VSS VDD _1348_ _1357_ core.pdc.row_out_n\[13\] _1336_ VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_135_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_45 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_100_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_153 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_85_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2920_ VSS VDD _0638_ _0708_ _0812_ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk2\[14\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[14\] core.ndc.rowon_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_90_498 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2851_ VDD VSS _0746_ core.cnb.shift_register_r\[9\] VSS VDD sky130_fd_sc_hd__inv_2
X_1802_ VDD VSS _1062_ core.ndc.col_out\[31\] _1126_ _1299_ _1251_ _1296_ VSS VDD
+ sky130_fd_sc_hd__a221o_4
X_2782_ VDD VSS _0678_ core.cnb.shift_register_r\[14\] VSS VDD sky130_fd_sc_hd__inv_2
X_1733_ VDD VSS core.ndc.col_out_n\[17\] _1258_ VSS VDD sky130_fd_sc_hd__buf_2
X_1664_ VSS VDD _1035_ _1198_ _1194_ _1075_ core.ndc.col_out_n\[9\] _1205_ VSS VDD
+ sky130_fd_sc_hd__o221a_2
XANTENNA__1934__B _1069_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_131_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1595_ VSS VDD _1045_ _1145_ _1079_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2111__A _1413_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2216_ VDD VSS _0239_ _0248_ _0243_ _0249_ VSS VDD sky130_fd_sc_hd__or3_1
X_3196_ VSS VDD net63 core.osr.next_sample_count_w\[4\] net77 core.osr.sample_count_r\[4\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2147_ VSS VDD core.cnb.average_counter_r\[1\] _0191_ core.cnb.average_counter_r\[0\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_93_281 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2078_ VSS VDD _0065_ _0095_ _0147_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2434__A1 core.pdc.rowoff_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2434__B2 _1325_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1945__A0 _1069_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout86_A net87 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1860__A net14 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_44_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_genblk2\[5\].buf_n_rowonn_A core.ndc.rowon_bottotop_n\[5\] VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_111_82 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk1\[29\].buf_n_coln VDD VSS core.ndc.col_out_n\[29\] nmatrix_col_core_n_buffered\[29\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_0_clk_dig_dummy_A cgen/clk_dig_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3050_ VSS VDD _0877_ _0894_ _0938_ VSS VDD sky130_fd_sc_hd__nand2b_1
XFILLER_96_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2585__B _1067_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2001_ VSS VDD _1162_ _1409_ _0094_ _1053_ VSS VDD sky130_fd_sc_hd__a21oi_2
XFILLER_90_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_284 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2903_ VDD VSS _0795_ _0784_ VSS VDD sky130_fd_sc_hd__inv_2
X_2834_ VSS VDD _0636_ _0728_ _0729_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__3103__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2765_ VSS VDD core.cnb.shift_register_r\[16\] _0638_ _0661_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2696_ VSS VDD _0519_ _0356_ _0528_ _0596_ VSS VDD sky130_fd_sc_hd__o21a_1
X_1716_ VSS VDD _1164_ _1127_ _1246_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1647_ VSS VDD _1190_ core.ndc.col_out_n\[8\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_116_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1578_ VSS VDD _1126_ _1129_ _1130_ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk1\[31\].buf_n_coln VDD VSS core.ndc.col_out_n\[31\] nmatrix_col_core_n_buffered\[31\]
+ VSS VDD sky130_fd_sc_hd__buf_6
X_3179_ VSS VDD net58 core.osr.next_result_w\[19\] net70 core.osr.result_r\[19\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_54_421 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_25_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2016__A core.pdc.col_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_373 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_248 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1590__A _1131_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_66_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_122_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3126__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1749__B _1177_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2550_ VSS VDD core.cnb.data_register_r\[0\] _0473_ _0474_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2481_ VSS VDD core.pdc.row_out_n\[14\] core.pdc.rowoff_out_n\[14\] core.pdc.rowon_out_n\[14\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_1501_ VSS VDD _1054_ _1061_ _1060_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1432_ VSS VDD _0992_ _0996_ _0995_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3102_ VDD VSS core.cnb.is_sampling_w net84 _0002_ clknet_2_0__leaf_clk_dig_dummy
+ VSS VDD sky130_fd_sc_hd__dfstp_1
Xgenblk2\[2\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[2\] core.pdc.row_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_83_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3033_ VSS VDD _0895_ _0920_ _0921_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_51_413 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_102_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1675__A _1138_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2817_ VDD VSS _0712_ _0711_ VSS VDD sky130_fd_sc_hd__inv_2
X_2748_ VSS VDD core.cnb.shift_register_r\[13\] _0644_ core.cnb.shift_register_r\[12\]
+ VSS VDD sky130_fd_sc_hd__nor2_2
X_2679_ VDD VSS _1008_ _0367_ _0524_ _0581_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_86_321 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_86_387 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2566__D _0482_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1842__A2 _1328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1981_ VDD VSS core.pdc.col_out_n\[5\] core.pdc.col_out\[5\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_61_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2602_ VSS VDD _0515_ core.cnb.result_out\[11\] _0438_ _0514_ VSS VDD sky130_fd_sc_hd__mux2_1
X_2533_ VSS VDD _0020_ _0458_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2464_ VSS VDD core.ndc.row_out_n\[11\] core.ndc.rowoff_out_n\[11\] core.ndc.rowon_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2395_ VDD VSS _0406_ _0405_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_3016_ VSS VDD _0902_ _0904_ _0903_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2086__A2 _1173_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[9\].buf_p_rowonn_A core.pdc.rowon_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_298 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_98_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2010__A2 _1395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2013__B _1101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1588__A1 _1137_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1762__B _1275_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2180_ VSS VDD _0208_ _0219_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1512__A1 _1069_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_74_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1579__A1 _1121_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1964_ VSS VDD _0065_ _0066_ _0067_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1579__B2 _1125_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1895_ VSS VDD _1305_ core.ndc.rowon_bottotop_n\[5\] _1308_ VSS VDD sky130_fd_sc_hd__nor2_2
X_2516_ VSS VDD _0012_ _0449_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2447_ VSS VDD _1374_ core.ndc.rowon_out_n\[8\] core.pdc.rowon_out_n\[15\] VSS VDD
+ sky130_fd_sc_hd__nand2_1
XFILLER_124_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2378_ VSS VDD core.osr.next_result_w\[19\] _0392_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_17_25 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2008__B _0098_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_33_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[1\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[1\] core.pdc.rowon_out_n\[1\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_3_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_109_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1863__A _1347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xcgen VDD comp/clk cgen/clk_dig_out net18 net25 net26 net27 net28 net29 net30 net31
+ net32 net33 net19 net20 net21 net22 net23 net3 net4 net5 net6 net7 net8 core.cnb.enable_loop_out
+ net24 decision_finish_comp_n net54 sample_nmatrix_cgen net55 sample_pmatrix_cgen
+ net35 VSS VSS adc_clkgen_with_edgedetect
XFILLER_87_471 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input29_A config_2_in[5] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_74_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_128_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_128_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1680_ VSS VDD _1217_ _1218_ _1152_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2301_ VDD VSS _0325_ _0324_ VSS VDD sky130_fd_sc_hd__inv_2
X_2232_ VSS VDD _0261_ _0263_ _0257_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2163_ VSS VDD _0205_ _0207_ _0206_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_80_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2094_ VDD VSS core.pdc.col_out_n\[23\] core.pdc.col_out\[23\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_62_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1667__B _1057_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2996_ VSS VDD _1113_ _0689_ _0886_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1947_ VSS VDD _1259_ _1399_ _1397_ _1224_ core.pdc.col_out_n\[1\] _1402_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
X_1878_ VSS VDD core.ndc.rowoff_out_n\[8\] _1314_ _1357_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1683__A _1220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_246 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3032__B _1104_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_411 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk2\[7\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[7\] core.pdc.row_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_90_433 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_455 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_90_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2850_ VSS VDD _0744_ _0731_ _0745_ _0725_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1801_ VSS VDD _1272_ _1084_ _1299_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2781_ VSS VDD _0666_ _0677_ _0676_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1732_ VSS VDD _1258_ _1257_ _1256_ _1255_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_116_126 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1663_ VSS VDD _1205_ _1110_ _1204_ VSS VDD sky130_fd_sc_hd__or2_1
X_1594_ VSS VDD _1074_ _1143_ _1144_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2111__B _1101_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2215_ VSS VDD _0246_ _0248_ _0247_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_85_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3195_ VSS VDD net63 core.osr.next_sample_count_w\[3\] net77 core.osr.sample_count_r\[3\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2146_ VDD VSS _0190_ core.cnb.average_counter_r\[3\] VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2682__A2 core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2077_ VDD VSS _0146_ _0111_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__3182__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1678__A core.ndc.col_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2979_ VSS VDD _0868_ _0870_ _0869_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_30_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1945__A1 _1067_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1860__B core.cnb.data_register_r\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[2\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[2\] core.pdc.col_out_n\[2\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1770__B _1095_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2000_ VDD VSS core.pdc.col_out_n\[7\] core.pdc.col_out\[7\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2902_ VSS VDD _0053_ _0794_ _0781_ _0793_ _1076_ _0688_ VSS VDD sky130_fd_sc_hd__a32o_1
X_2833_ VSS VDD _0668_ _0728_ _0637_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_77_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2764_ VSS VDD _0646_ _0660_ _0659_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1715_ VDD VSS core.ndc.col_out\[14\] core.ndc.col_out_n\[14\] VSS VDD sky130_fd_sc_hd__inv_2
X_2695_ VSS VDD _0593_ _0594_ _0045_ _0595_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1646_ VSS VDD _1190_ _1189_ _1185_ _1181_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__2122__A _1396_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1577_ VSS VDD _1128_ _1127_ _1129_ _1082_ VSS VDD sky130_fd_sc_hd__a21oi_2
Xgenblk2\[4\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[4\] core.ndc.row_out_n\[4\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1680__B _1152_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3178_ VSS VDD net58 core.osr.next_result_w\[18\] net69 core.osr.result_r\[18\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2129_ VDD VSS _1126_ _1393_ core.pdc.col_out\[31\] _1121_ _1391_ _0175_ VSS VDD
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_25_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3099__S _0241_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_41_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input11_A config_1_in[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_60 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2207__A _0240_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2582__A1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2480_ VSS VDD core.pdc.rowon_out_n\[13\] core.pdc.rowoff_out_n\[13\] core.pdc.row_out_n\[13\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_56_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2582__B2 _1104_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1500_ VSS VDD _1059_ _1060_ _1057_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1431_ VSS VDD _0993_ _0994_ _0995_ VSS VDD sky130_fd_sc_hd__nor2_1
X_3101_ VSS VDD clknet_2_0__leaf_clk_dig_dummy core.cnb.next_conv_finished_w net84
+ net37 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_55_219 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3032_ VSS VDD _0917_ _1104_ _0920_ _0919_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_83_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_425 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2816_ VSS VDD _0710_ _0711_ _0664_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1956__A core.pdc.col_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1675__B _1177_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2747_ VSS VDD _0641_ _0643_ _0642_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2678_ VSS VDD _0578_ _0579_ _0043_ _0580_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1629_ VSS VDD _1085_ _1043_ _1118_ _1175_ VSS VDD sky130_fd_sc_hd__o21a_1
XANTENNA_input3_A config_1_in[10] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_300 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_117_71 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_cgen_ena_in core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_358 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_93_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1980_ VSS VDD _1259_ _0076_ _0074_ _1224_ core.pdc.col_out_n\[5\] _0078_ VSS VDD
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1776__A _1033_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2601_ VDD VSS _1309_ _0514_ _0513_ VSS VDD sky130_fd_sc_hd__xor2_1
X_2532_ VSS VDD _0458_ net9 net54 core.cnb.sampled_avg_control_r\[1\] VSS VDD sky130_fd_sc_hd__mux2_1
X_2463_ VSS VDD core.ndc.row_out_n\[10\] core.ndc.rowoff_out_n\[10\] core.ndc.rowon_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2394_ VSS VDD _0403_ _0404_ _0405_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_56_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3015_ VSS VDD _0901_ _0903_ _1312_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_325 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_380 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk1\[8\].buf_n_coln_A core.ndc.col_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2010__A3 _1085_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3116__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_fanout61_A net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_112 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[13\].buf_p_rown_A core.pdc.row_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_155 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1963_ VSS VDD _0066_ _1170_ _1400_ _1145_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1894_ VSS VDD core.pdc.rowon_out_n\[2\] _1366_ _1368_ VSS VDD sky130_fd_sc_hd__nand2_2
XANTENNA__1579__A2 _1124_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2528__A1 net54 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3139__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2515_ VSS VDD _0449_ core.cnb.shift_register_r\[11\] _0444_ core.cnb.shift_register_r\[10\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_2446_ VSS VDD core.ndc.rowon_out_n\[7\] _0429_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2130__A core.pdc.col_out\[31\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2377_ VSS VDD _0392_ _0391_ _0240_ _0390_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_68_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk1\[7\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[7\] core.pdc.col_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_137_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_58_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2694__B core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2455__B1 core.pdc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_23_91 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_99_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2300_ VDD VSS _0315_ _0306_ _0314_ _0324_ VSS VDD sky130_fd_sc_hd__a21oi_1
X_2231_ VDD VSS _0252_ core.cnb.result_out\[2\] _0262_ core.osr.next_result_w\[2\]
+ VSS VDD sky130_fd_sc_hd__a21o_1
X_2162_ VSS VDD core.cnb.shift_register_r\[4\] core.cnb.shift_register_r\[5\] _0206_
+ VSS VDD sky130_fd_sc_hd__nor2_1
Xgenblk2\[9\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[9\] core.ndc.row_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2093_ VSS VDD core.pdc.col_out_n\[23\] _0155_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_80_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__3189__RESET_B net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2995_ VSS VDD _0883_ _0885_ _0879_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_119_135 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3118__RESET_B net86 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1946_ VSS VDD _1401_ _1402_ _1155_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1877_ VSS VDD _1356_ core.pdc.row_out_n\[12\] _1354_ VSS VDD sky130_fd_sc_hd__nor2_2
XANTENNA__1964__A _0065_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2429_ VSS VDD _1342_ _1314_ _0426_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_28_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2019__B _1135_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1858__B core.ndc.rowoff_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_100_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_69_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xgenblk1\[4\].buf_n_coln VDD VSS core.ndc.col_out_n\[4\] nmatrix_col_core_n_buffered\[4\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_62_114 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_85_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_309 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1768__B _1279_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1651__A1 _1077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1800_ VDD VSS core.ndc.col_out\[30\] core.ndc.col_out_n\[30\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_86_6 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2780_ VDD VSS _0676_ _0675_ VSS VDD sky130_fd_sc_hd__inv_2
X_1731_ VSS VDD _1165_ _1257_ _1188_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1662_ VSS VDD _1043_ _1203_ _1204_ _1199_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1593_ VSS VDD _1142_ _1103_ _1143_ _1141_ VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_85_206 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_3194_ VSS VDD net62 core.osr.next_sample_count_w\[2\] net75 core.osr.sample_count_r\[2\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2214_ VSS VDD core.cnb.result_out\[1\] _0247_ core.osr.result_r\[1\] VSS VDD sky130_fd_sc_hd__nand2_1
X_2145_ VDD VSS _0179_ _0188_ _0189_ _0185_ VSS VDD sky130_fd_sc_hd__o21bai_1
XFILLER_53_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2076_ VDD VSS core.pdc.col_out_n\[19\] core.pdc.col_out\[19\] VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_53_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2978_ VSS VDD _0865_ _0866_ _0869_ _1114_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1929_ VSS VDD _1387_ core.pdc.rowon_out_n\[15\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1694__A _1105_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_130_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1869__A net14 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_88 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1936__A2 _1284_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_130 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2649__B1 _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_220 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1779__A core.ndc.col_out\[25\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3074__B1 _1312_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_253 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2901_ VSS VDD _0792_ _0794_ _0791_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2832_ VDD VSS _0727_ _0726_ VSS VDD sky130_fd_sc_hd__inv_2
X_2763_ VSS VDD _0659_ _0650_ _0641_ VSS VDD sky130_fd_sc_hd__nand2_2
X_1714_ VDD VSS core.ndc.col_out_n\[14\] _1245_ VSS VDD sky130_fd_sc_hd__buf_2
X_2694_ VSS VDD _0542_ _0595_ core.cnb.result_out\[7\] VSS VDD sky130_fd_sc_hd__nand2_1
X_1645_ VSS VDD _1187_ _1189_ _1188_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2122__B _1188_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1576_ VSS VDD _1057_ _1128_ _1087_ VSS VDD sky130_fd_sc_hd__nor2_2
Xgenblk2\[10\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[10\] core.ndc.rowon_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1961__B _1088_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3177_ VSS VDD net57 core.osr.next_result_w\[17\] net69 core.osr.result_r\[17\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__2792__B _0208_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2128_ VDD VSS _0175_ _1401_ _1092_ VSS VDD sky130_fd_sc_hd__and2_1
X_2059_ VSS VDD core.pdc.col_out_n\[15\] _0137_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_41_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2967__B _1076_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_122_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_122_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1599__A _1148_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2582__A2 _0439_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1430_ VSS VDD core.osr.osr_mode_r\[2\] _0990_ _0994_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__3172__CLK net58 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3100_ VSS VDD _0064_ _0981_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_3031_ VSS VDD _0918_ _0919_ _0916_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_51_437 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2117__B _1235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2815_ VSS VDD _0709_ _0660_ _0710_ _0661_ VSS VDD sky130_fd_sc_hd__nand3_1
XANTENNA__2133__A core.cnb.sampled_avg_control_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2746_ VDD VSS _0642_ core.cnb.shift_register_r\[16\] VSS VDD sky130_fd_sc_hd__inv_2
X_2677_ VSS VDD core.osr.next_result_w\[5\] _0580_ _0542_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1972__A _0065_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1781__B1 _1035_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1628_ VSS VDD _1172_ _1174_ _1173_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1559_ VDD VSS _1113_ core.cnb.data_register_r\[6\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_86_367 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_14_128 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_77_21 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2600_ VSS VDD _1328_ _0501_ _0513_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2531_ VSS VDD _0019_ _0457_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2462_ VSS VDD core.ndc.row_out_n\[9\] core.ndc.rowoff_out_n\[9\] core.ndc.rowon_out_n\[9\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2393_ VDD VSS _0404_ _0401_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3014_ VSS VDD _0902_ _1312_ _0901_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_83_337 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2729_ VSS VDD _0624_ _0626_ _0625_ VSS VDD sky130_fd_sc_hd__nand2_1
Xgenblk2\[7\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[7\] core.ndc.rowon_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2310__B _0255_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_fanout54_A net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[9\].buf_n_coln VDD VSS core.ndc.col_out_n\[9\] nmatrix_col_core_n_buffered\[9\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_137_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_71 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_167 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1962_ VSS VDD _1110_ _0065_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1893_ VDD VSS _1368_ _1367_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1984__A0 _1118_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2514_ VSS VDD _0011_ _0448_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2445_ VSS VDD _0429_ _1351_ _1364_ VSS VDD sky130_fd_sc_hd__or2_1
X_2376_ VSS VDD _0391_ core.osr.result_r\[18\] core.osr.result_r\[19\] _0384_ VSS
+ VDD sky130_fd_sc_hd__nand3b_1
XFILLER_56_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_137_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_58_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_47_337 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_114_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_139_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2230_ VSS VDD _0262_ _0261_ _0260_ _0255_ VSS VDD sky130_fd_sc_hd__and3_1
X_2161_ VSS VDD core.cnb.shift_register_r\[2\] core.cnb.shift_register_r\[3\] _0205_
+ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_93_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_65_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2092_ VSS VDD _0155_ _0154_ _0153_ _0152_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_0_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2994_ VSS VDD _0884_ _0879_ _0883_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__3106__CLK clknet_2_2__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1945_ VSS VDD _1401_ _1067_ _1400_ _1069_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_119_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1876_ VSS VDD _1311_ _1355_ _1356_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2428_ VSS VDD _1334_ _1315_ core.ndc.row_out_n\[9\] VSS VDD sky130_fd_sc_hd__nor2_1
X_2359_ VDD VSS _0373_ _0377_ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_56_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_351 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_13 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_100_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_60_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2051__A _1396_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input34_A rst_n VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_281 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_178 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3129__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1730_ VSS VDD _1100_ _1256_ _1213_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1661_ VSS VDD _1043_ _1203_ _1202_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1592_ VSS VDD _1103_ _1142_ _1112_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3193_ VSS VDD net62 core.osr.next_sample_count_w\[1\] net75 core.osr.sample_count_r\[1\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2213_ VSS VDD _0244_ _0246_ _0245_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2144_ VDD VSS _0188_ _0187_ VSS VDD sky130_fd_sc_hd__inv_2
X_2075_ VSS VDD core.pdc.col_out_n\[19\] _0145_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_53_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2136__A core.cnb.sampled_avg_control_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2977_ VSS VDD _0867_ _0868_ _1087_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1928_ VSS VDD _1387_ _1038_ _1030_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_30_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1859_ VSS VDD _1325_ _1318_ _1344_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_122_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_115_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2658__A1 core.osr.next_result_w\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_44_126 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3083__A1 _0758_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2649__A1 core.osr.next_result_w\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_232 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_265 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2900_ VSS VDD _0793_ _0791_ _0792_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1795__A _1272_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2831_ VSS VDD _0725_ _0723_ _0726_ _0724_ VSS VDD sky130_fd_sc_hd__nand3_2
X_2762_ VSS VDD _0206_ _0657_ _0658_ core.cnb.shift_register_r\[7\] VSS VDD sky130_fd_sc_hd__nand3_1
X_1713_ VSS VDD _1245_ _1244_ _1241_ _1239_ VSS VDD sky130_fd_sc_hd__and3_1
X_2693_ VSS VDD _0395_ _0594_ net40 VSS VDD sky130_fd_sc_hd__nand2_1
X_1644_ VDD VSS _1188_ _1032_ VSS VDD sky130_fd_sc_hd__buf_2
X_1575_ VSS VDD _1053_ _1042_ _1127_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_112_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3176_ VSS VDD net56 core.osr.next_result_w\[16\] net68 core.osr.result_r\[16\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_26_115 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2127_ VDD VSS core.pdc.col_out_n\[30\] core.pdc.col_out\[30\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2058_ VSS VDD _0137_ _0136_ _0132_ _0130_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__3173__RESET_B net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A net85 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[15\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[15\] core.pdc.rowon_out_n\[15\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_106_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1854__A2 _1340_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3056__A1 _1312_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_99 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_31_92 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3030_ VDD VSS _0918_ _0847_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_31_140 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2814_ VSS VDD _0706_ _0709_ _0708_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_82_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2745_ VSS VDD core.cnb.shift_register_r\[10\] core.cnb.shift_register_r\[11\] _0641_
+ VSS VDD sky130_fd_sc_hd__nor2_1
X_2676_ VSS VDD _0395_ _0579_ net53 VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1781__A1 _1259_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1627_ VSS VDD _1032_ _1173_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1972__B _0072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1558_ VDD VSS _1112_ _1111_ VSS VDD sky130_fd_sc_hd__inv_2
X_1489_ VSS VDD _1037_ _1048_ _1049_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_86_379 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3159_ VSS VDD net62 _0049_ net74 net44 VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__2043__B _1163_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_117_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2530_ VSS VDD _0457_ net2 net54 core.cnb.sampled_avg_control_r\[0\] VSS VDD sky130_fd_sc_hd__mux2_1
X_2461_ VSS VDD core.ndc.row_out_n\[7\] core.ndc.rowoff_out_n\[7\] core.ndc.rowon_out_n\[7\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2392_ VDD VSS _0403_ core.osr.sample_count_r\[3\] VSS VDD sky130_fd_sc_hd__inv_2
X_3013_ VSS VDD _0697_ _0900_ _0901_ _0847_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_83_349 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2128__B _1092_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2728_ VSS VDD core.osr.next_result_w\[15\] _0625_ _0568_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2659_ VDD VSS _0564_ _0563_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2703__B1 core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_154 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_68_891 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2038__B _1095_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_128_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_74_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1961_ VSS VDD _1413_ _1412_ _1088_ VSS VDD sky130_fd_sc_hd__nand2_2
X_1892_ VSS VDD _1362_ _1029_ _1367_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1984__A1 _1112_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2513_ VSS VDD _0448_ core.cnb.shift_register_r\[10\] _0444_ core.cnb.shift_register_r\[9\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_2444_ VDD VSS core.ndc.rowon_out_n\[6\] _0428_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_124_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2375_ VSS VDD _0390_ _0383_ core.osr.result_r\[18\] _0377_ core.osr.result_r\[19\]
+ VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_56_305 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_500 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_65_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__3185__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1672__B1 _1206_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1975__A1 _1141_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_55 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_128_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_99_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_99_86 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk_dig_dummy VSS VDD cgen/clk_dig_out clknet_0_clk_dig_dummy VSS VDD sky130_fd_sc_hd__clkbuf_16
X_2160_ VDD VSS _0204_ _0203_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_17_5 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2091_ VSS VDD _0096_ _0154_ _1101_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_93_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_93_477 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_382 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1798__A _1272_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2993_ VSS VDD _0882_ _0883_ _0868_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_9_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1944_ VSS VDD _1388_ _1400_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1875_ VDD VSS _1355_ _1024_ VSS VDD sky130_fd_sc_hd__inv_2
X_2427_ VSS VDD _1337_ core.ndc.row_out_n\[8\] core.pdc.rowoff_out_n\[0\] VSS VDD
+ sky130_fd_sc_hd__nand2_1
XFILLER_88_238 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2358_ VDD VSS core.osr.next_result_w\[15\] _0376_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_56_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2289_ VSS VDD core.osr.result_r\[9\] core.cnb.result_out\[9\] _0314_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_60_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__2051__B _1152_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_125_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input27_A config_2_in[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_293 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__2242__A core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1660_ VDD VSS _1202_ _1201_ VSS VDD sky130_fd_sc_hd__inv_2
X_1591_ VDD VSS _1104_ _1105_ _1088_ _1141_ VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_124_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2896__B _1076_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3192_ VDD VSS core.osr.sample_count_r\[0\] net74 core.osr.next_sample_count_w\[0\]
+ net62 VSS VDD sky130_fd_sc_hd__dfstp_1
X_2212_ VDD VSS _0245_ core.osr.result_r\[1\] VSS VDD sky130_fd_sc_hd__inv_2
X_2143_ VSS VDD _0176_ _0186_ _0187_ core.cnb.sampled_avg_control_r\[2\] VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_93_230 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_93_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2074_ VSS VDD _0145_ _0144_ _0143_ _0142_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_14_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2976_ VSS VDD _0865_ _0867_ _0866_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1927_ VSS VDD core.pdc.rowon_out_n\[14\] core.ndc.rowon_out_n\[0\] _1386_ VSS VDD
+ sky130_fd_sc_hd__nand2_2
XFILLER_30_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1858_ VSS VDD _1343_ core.pdc.row_out_n\[8\] core.ndc.rowoff_out_n\[0\] VSS VDD
+ sky130_fd_sc_hd__nand2_1
X_1789_ VDD VSS core.ndc.col_out_n\[27\] core.ndc.col_out\[27\] VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1991__A core.pdc.col_out_n\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_130_110 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1885__B core.ndc.rowon_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_29_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_244 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk2\[10\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[10\] core.pdc.row_out_n\[10\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2830_ VDD VSS _0725_ _0649_ VSS VDD sky130_fd_sc_hd__buf_2
X_2761_ VDD VSS _0657_ core.cnb.shift_register_r\[6\] VSS VDD sky130_fd_sc_hd__inv_2
X_2692_ VDD VSS _0588_ _0592_ _0593_ _0591_ VSS VDD sky130_fd_sc_hd__o21bai_1
X_1712_ VSS VDD _1244_ _1034_ _1243_ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_6_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1643_ VSS VDD _1186_ _1113_ _1187_ _1043_ VSS VDD sky130_fd_sc_hd__o21ai_2
X_1574_ VDD VSS _1126_ _1110_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_86_506 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_110 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_3175_ VSS VDD net58 core.osr.next_result_w\[15\] net70 core.osr.result_r\[15\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_26_127 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2126_ VSS VDD core.pdc.col_out_n\[30\] _0174_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_54_447 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2057_ VSS VDD _0136_ _1034_ _0135_ VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1986__A _1206_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2959_ VSS VDD _0776_ _0791_ _0851_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__3142__RESET_B net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3119__CLK clknet_2_0__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_106_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2057__A _1034_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_40_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2813_ VSS VDD _0707_ _0708_ _0206_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2007__A0 _1161_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2744_ VDD VSS _0639_ _0640_ VSS VDD sky130_fd_sc_hd__buf_6
X_2675_ VDD VSS _0573_ _0577_ _0578_ _0576_ VSS VDD sky130_fd_sc_hd__o21bai_1
XANTENNA__1781__A2 _1220_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1626_ VDD VSS _1172_ _1171_ VSS VDD sky130_fd_sc_hd__inv_2
X_1557_ VSS VDD _1085_ _1065_ _1111_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_98_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1488_ VSS VDD _1043_ _1048_ _1047_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3158_ VSS VDD net60 _0048_ net74 net43 VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_36_49 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2109_ VDD VSS _0161_ _0162_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_3089_ VSS VDD _0966_ _0973_ _0974_ _0969_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_22_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2978__C _1114_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_genblk2\[2\].buf_n_rown_A core.ndc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1565__S _1077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2460_ VSS VDD core.ndc.row_out_n\[6\] core.ndc.rowoff_out_n\[6\] core.ndc.rowon_out_n\[6\]
+ VSS VDD sky130_fd_sc_hd__nand2_1
X_2391_ VDD VSS core.osr.next_sample_count_w\[2\] _0402_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_en_bit_n[2] core.cnb.pswitch_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3012_ VSS VDD _0799_ _0900_ _0697_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_51_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_225 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2727_ VSS VDD core.osr.next_result_w\[17\] _0624_ _1002_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1983__B _1279_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2658_ VDD VSS _0393_ core.osr.next_result_w\[3\] _0562_ _0563_ net51 VSS VDD sky130_fd_sc_hd__a22o_1
X_1609_ VSS VDD _1076_ _1156_ _1145_ _1157_ VSS VDD sky130_fd_sc_hd__o21a_1
X_2589_ VSS VDD _0503_ _0505_ _0504_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_47_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input1_A clk_vcm VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_103_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[11\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[11\] core.pdc.col_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_88_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_37_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1960_ VSS VDD _1409_ _1412_ _1036_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_53_91 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1891_ VDD VSS _1366_ _1365_ VSS VDD sky130_fd_sc_hd__inv_2
X_2512_ VSS VDD _0010_ _0447_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_52_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2443_ VSS VDD _1379_ _0428_ _1368_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2374_ VSS VDD core.osr.next_result_w\[18\] _0389_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_83_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_512 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_137_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_137_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_genblk1\[19\].buf_n_coln_A core.ndc.col_out_n\[19\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_497 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_361 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xgenblk2\[3\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[3\] core.ndc.rowon_out_n\[3\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__2065__A _0065_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_130_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xgenblk2\[15\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[15\] core.pdc.row_out_n\[15\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_90_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_23_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2090_ VSS VDD _0139_ _0153_ _1235_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_93_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_350 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_361 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_93_489 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2992_ VSS VDD _0863_ _0882_ _0881_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_9_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_genblk1\[9\].buf_p_coln_A core.pdc.col_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1943_ VDD VSS _1399_ _1398_ VSS VDD sky130_fd_sc_hd__inv_2
X_1874_ VSS VDD core.ndc.rowoff_out_n\[8\] _1349_ _1354_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1753__S _1034_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_206 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2426_ VSS VDD _1343_ core.ndc.row_out_n\[7\] _1361_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_88_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2357_ VSS VDD _0369_ _0376_ _0375_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2288_ VDD VSS _0313_ core.osr.next_result_w\[8\] _0252_ _0312_ VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_84_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3167__RESET_B net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_44_49 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1501__B _1060_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_100_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_109_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_125_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1899__A _1371_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_404 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__3175__CLK net58 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1590_ VSS VDD _1131_ _1139_ _1140_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2211_ VDD VSS _0244_ core.cnb.result_out\[1\] VSS VDD sky130_fd_sc_hd__inv_2
X_3191_ VDD VSS core.cnb.data_register_r\[11\] net82 _0061_ clknet_2_1__leaf_clk_dig_dummy
+ VSS VDD sky130_fd_sc_hd__dfstp_2
X_2142_ VDD VSS _0186_ core.cnb.sampled_avg_control_r\[0\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_38_114 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_2073_ VSS VDD _0144_ _1033_ _0113_ VSS VDD sky130_fd_sc_hd__or2_1
Xgenblk2\[12\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[12\] core.ndc.row_out_n\[12\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_46_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2975_ VSS VDD _0795_ _0866_ _0864_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1926_ VSS VDD _1385_ _1386_ _1027_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_30_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1857_ VDD VSS _1342_ _1024_ _1336_ _1343_ VSS VDD sky130_fd_sc_hd__a21o_1
X_1788_ VSS VDD core.ndc.col_out_n\[27\] _1293_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_130_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_39_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2409_ VSS VDD _0414_ _0417_ core.osr.sample_count_r\[6\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_44_106 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_106_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_401 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_434 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_29_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1609__A1 _1076_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2253__A core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2760_ VSS VDD _0648_ _0656_ _0655_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2691_ VSS VDD core.osr.next_result_w\[9\] _1019_ _0592_ _0537_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1711_ VSS VDD _1243_ _1202_ _1054_ _1242_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__3068__B _0799_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1642_ VSS VDD _1116_ _1186_ _1117_ VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_6_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1573_ VSS VDD _1095_ _1125_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__3084__A _1022_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_518 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3174_ VSS VDD net58 core.osr.next_result_w\[14\] net70 core.osr.result_r\[14\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2125_ VSS VDD _0174_ _0173_ _0171_ _0170_ VSS VDD sky130_fd_sc_hd__and3_1
X_2056_ VSS VDD _1242_ _0134_ _0135_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_41_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2958_ VSS VDD _0849_ _0850_ _0755_ VSS VDD sky130_fd_sc_hd__nand2_1
Xgenblk1\[16\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[16\] core.pdc.col_out_n\[16\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1909_ VSS VDD _1340_ core.pdc.rowon_out_n\[7\] core.pdc.rowoff_out_n\[8\] VSS VDD
+ sky130_fd_sc_hd__nand2_1
X_2889_ VSS VDD _0052_ _0782_ _0781_ _0780_ _0482_ _0758_ VSS VDD sky130_fd_sc_hd__a32o_1
XFILLER_103_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3182__RESET_B net86 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_122_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_15_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2073__A _1033_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1417__A core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput50 VDD VSS result_out[6] net50 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_48_286 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2812_ VSS VDD core.cnb.shift_register_r\[7\] _0657_ _0707_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_72_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2007__A1 _1229_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2743_ VSS VDD _0636_ _0638_ _0639_ VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_68_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2674_ VSS VDD core.osr.next_result_w\[7\] _1019_ _0577_ _0537_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1625_ VSS VDD _1156_ _1171_ _1170_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1556_ VDD VSS _1110_ _1039_ VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1487_ VSS VDD _1046_ _1047_ _1044_ VSS VDD sky130_fd_sc_hd__nor2_2
X_3157_ VSS VDD net59 _0047_ net72 net42 VSS VDD sky130_fd_sc_hd__dfrtp_1
X_2108_ VSS VDD _1131_ _0091_ _0161_ VSS VDD sky130_fd_sc_hd__nor2_1
X_3088_ VDD VSS _0973_ _0971_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1997__A _0091_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2039_ VSS VDD _0122_ _0121_ _0119_ _0117_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_52_16 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_462 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_77_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_92_329 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1700__A _1034_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[13\].buf_n_coln VDD VSS core.ndc.col_out_n\[13\] nmatrix_col_core_n_buffered\[13\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_9_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1996__B1 _1045_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[11\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[11\] core.pdc.rowon_out_n\[11\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_3_21 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2390_ VDD VSS _0401_ core.osr.is_last_sample _0400_ _0402_ VSS VDD sky130_fd_sc_hd__or3_1
XANTENNA_nmat_en_bit_n[1] core.cnb.pswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__3081__B _0691_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_3011_ VSS VDD _0689_ _0899_ _0057_ _1053_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_91_351 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__3109__CLK clknet_2_3__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[7\].buf_p_rown_A core.pdc.row_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2726_ VSS VDD core.osr.next_result_w\[19\] _0623_ _0533_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2441__A core.pdc.rowon_bottotop_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2657_ VSS VDD _0983_ _0562_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1608_ VSS VDD _1043_ _1156_ _1045_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2588_ VSS VDD _0501_ _0504_ _1300_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1539_ VSS VDD _1072_ _1095_ VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_103_11 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_103_66 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1520__A _1077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_128_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_88_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1890_ VSS VDD _1338_ _1028_ _1365_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2261__A core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2511_ VSS VDD _0447_ core.cnb.shift_register_r\[9\] _0444_ core.cnb.shift_register_r\[8\]
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_2442_ VSS VDD core.ndc.rowoff_out_n\[5\] core.ndc.rowon_out_n\[4\] _1311_ VSS VDD
+ sky130_fd_sc_hd__nand2_1
X_2373_ VSS VDD _0389_ _0240_ _0388_ _0387_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_83_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_524 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_181 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2709_ VSS VDD _0363_ _1011_ _0608_ _0518_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1515__A _1072_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_74_115 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_74_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_135_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_395 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2991_ VDD VSS _0881_ _0880_ VSS VDD sky130_fd_sc_hd__inv_2
X_1942_ VSS VDD _1398_ _1098_ _1394_ _1067_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1873_ VDD VSS core.pdc.row_out_n\[11\] _1353_ VSS VDD sky130_fd_sc_hd__inv_2
Xgenblk2\[8\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[8\] core.pdc.rowon_out_n\[8\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_134_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2425_ VDD VSS core.ndc.row_out_n\[6\] _0425_ VSS VDD sky130_fd_sc_hd__inv_2
X_2356_ VDD VSS _0375_ _0374_ VSS VDD sky130_fd_sc_hd__inv_2
X_2287_ VSS VDD _0252_ _0313_ core.cnb.result_out\[8\] VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_71_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_32 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2530__A0 core.cnb.sampled_avg_control_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_262 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xgenblk1\[23\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[23\] core.pdc.col_out_n\[23\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_18_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_109_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_genblk1\[0\].buf_n_coln_A core.ndc.col_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2210_ VDD VSS _0243_ core.osr.result_r\[0\] VSS VDD sky130_fd_sc_hd__inv_2
X_3190_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0060_ net81 core.cnb.data_register_r\[10\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
X_2141_ VDD VSS _0184_ _0183_ _0177_ _0185_ VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_38_126 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_265 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2072_ VSS VDD _0084_ _0143_ _1275_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2974_ VDD VSS _0472_ _0783_ _0864_ _0865_ VSS VDD sky130_fd_sc_hd__a21o_1
X_1925_ VSS VDD _1029_ _1385_ _1023_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1856_ VDD VSS _1342_ _1301_ VSS VDD sky130_fd_sc_hd__buf_2
X_1787_ VSS VDD _1293_ _1292_ _1291_ _1290_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_115_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_89_505 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_130_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2408_ VSS VDD core.osr.sample_count_r\[6\] _0414_ _0416_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2339_ VDD VSS _0360_ _0359_ _0271_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_29_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_111_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2579__B1 core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[18\].buf_n_coln VDD VSS core.ndc.col_out_n\[18\] nmatrix_col_core_n_buffered\[18\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_20_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_106_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_136_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_136_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1857__A2 _1342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input32_A config_2_in[8] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3142__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2690_ VSS VDD _0589_ _0591_ _0590_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_61_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1710_ VSS VDD _1060_ _1242_ _1117_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1641_ VDD VSS _1184_ _1185_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_6_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1572_ VSS VDD _1124_ _1068_ _1078_ _1123_ VSS VDD sky130_fd_sc_hd__o21a_2
XFILLER_112_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xgenblk1\[20\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[20\] core.ndc.col_out_n\[20\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_3173_ VSS VDD net61 core.osr.next_result_w\[13\] net73 core.osr.result_r\[13\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__1613__A core.ndc.col_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2124_ VDD VSS _0172_ _0173_ VSS VDD sky130_fd_sc_hd__clkinv_2
X_2055_ VDD VSS _0134_ _0133_ VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__2444__A _0428_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2957_ VSS VDD _0846_ core.cnb.data_register_r\[1\] _0849_ _0848_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2888_ VSS VDD _0779_ _0782_ _0777_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1908_ VSS VDD core.pdc.rowon_out_n\[6\] _1377_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1839_ VDD VSS _1327_ _1328_ VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_103_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_103_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_2_3__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_3__leaf_clk_dig_dummy
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
XFILLER_66_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__2073__B _0113_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput51 VDD VSS result_out[7] net51 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput40 VDD VSS result_out[11] net40 VSS VDD sky130_fd_sc_hd__buf_2
X_2811_ VSS VDD _0635_ core.cnb.shift_register_r\[4\] _0706_ _0705_ VSS VDD sky130_fd_sc_hd__nand3_1
X_2742_ VSS VDD _0638_ _0205_ _0637_ VSS VDD sky130_fd_sc_hd__nand2_2
X_2673_ VSS VDD _0574_ _0576_ _0575_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1624_ VSS VDD _1169_ _1170_ _1045_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1555_ VSS VDD _1088_ _1037_ _1109_ _1103_ VSS VDD sky130_fd_sc_hd__o21ai_2
X_1486_ VDD VSS _1046_ _1045_ VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_100_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3156_ VSS VDD net59 _0046_ net71 net41 VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__3188__CLK clknet_2_1__leaf_clk_dig_dummy VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_3087_ VSS VDD _0970_ _0972_ _0971_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2107_ VDD VSS core.pdc.col_out\[27\] core.pdc.col_out_n\[27\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2038_ VSS VDD _0120_ _0121_ _1095_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_fanout82_A net83 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_77_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_133_31 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2068__B _1155_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2084__A _1039_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_en_bit_n[0] core.cnb.pswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_3010_ VSS VDD _0897_ _0781_ _0899_ _0898_ VSS VDD sky130_fd_sc_hd__nand3_1
XFILLER_77_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_363 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_2725_ VSS VDD _0616_ _0048_ _0622_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2656_ VSS VDD _0559_ _0540_ _0561_ _0560_ VSS VDD sky130_fd_sc_hd__nand3_1
X_1607_ VDD VSS _1155_ _1101_ VSS VDD sky130_fd_sc_hd__buf_2
X_2587_ VDD VSS _0503_ _0502_ VSS VDD sky130_fd_sc_hd__inv_2
X_1538_ VDD VSS core.ndc.col_out\[1\] core.ndc.col_out_n\[1\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_86_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1469_ VDD VSS _1031_ net14 VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_68_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_179 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_3139_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0029_ net79 core.cnb.result_out\[7\]
+ VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_103_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1801__A _1272_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[28\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[28\] core.pdc.col_out_n\[28\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_103_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_103_89 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_128_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xgenblk1\[30\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[30\] core.pdc.col_out_n\[30\]
+ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2510_ VSS VDD _0009_ _0446_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_2441_ VSS VDD _1382_ core.ndc.rowon_out_n\[3\] core.pdc.rowon_bottotop_n\[5\] VSS
+ VDD sky130_fd_sc_hd__nor2_2
X_2372_ VDD VSS _0383_ _0377_ core.osr.result_r\[18\] _0388_ VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__2449__A2 core.pdc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_116 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1621__A _1131_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_193 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2708_ VSS VDD _0606_ _0607_ _0519_ VSS VDD sky130_fd_sc_hd__nand2_1
X_2639_ VSS VDD _0518_ _0288_ _0537_ _0546_ VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_59_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_477 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2627__A _1002_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1531__A _1088_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2612__A2 _0395_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_128_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_139_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__2081__B _1284_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1706__A _1227_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_rowoff_n[5] core.ndc.rowoff_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[25\].buf_n_coln VDD VSS core.ndc.col_out_n\[25\] nmatrix_col_core_n_buffered\[25\]
+ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_48_60 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2990_ VSS VDD _0802_ _0880_ _0869_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1941_ VDD VSS _1397_ _1396_ VSS VDD sky130_fd_sc_hd__inv_2
X_1872_ VDD VSS _1353_ _1350_ _1352_ VSS VDD sky130_fd_sc_hd__or2_2
XFILLER_43_1 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2424_ VSS VDD _0425_ _1360_ _1346_ VSS VDD sky130_fd_sc_hd__or2_1
X_2355_ VSS VDD _0374_ _0251_ _0373_ VSS VDD sky130_fd_sc_hd__or2_1
X_2286_ VSS VDD _0310_ _0312_ _0311_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_44_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_109_11 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__3163__D core.osr.next_result_w\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_171 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk1\[15\].buf_n_coln_A core.ndc.col_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_34_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1572__A2 _1078_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2140_ VDD VSS _0184_ core.cnb.average_counter_r\[2\] VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_38_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2071_ VSS VDD _0081_ _0142_ _1213_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_93_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_182 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_93_299 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_2973_ VSS VDD _0864_ _0697_ _0655_ _0764_ VSS VDD sky130_fd_sc_hd__nand3b_1
X_1924_ VSS VDD _1384_ core.pdc.rowon_out_n\[13\] _1364_ VSS VDD sky130_fd_sc_hd__nor2_2
X_1855_ VSS VDD core.pdc.row_out_n\[7\] _1337_ _1341_ VSS VDD sky130_fd_sc_hd__nand2_2
X_1786_ VSS VDD _1106_ _1292_ _1188_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_89_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[2\].buf_p_rowonn_A core.pdc.rowon_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2407_ VDD VSS _0415_ core.osr.next_sample_count_w\[5\] VSS VDD sky130_fd_sc_hd__clkinv_2
X_2338_ VSS VDD _0353_ _0359_ _0358_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__2177__A _0210_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_2269_ VSS VDD _0296_ core.osr.next_result_w\[6\] VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__2276__B1 _0255_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[9] nmatrix_col_core_n_buffered\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[3\].buf_n_rowonn_A core.ndc.rowon_out_n\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_136_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_64 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_96_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_136_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input25_A config_2_in[1] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1640_ VSS VDD _1039_ _1183_ _1184_ VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__2550__A core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1571_ VSS VDD _1122_ _1123_ _1051_ VSS VDD sky130_fd_sc_hd__nand2_1
X_3172_ VSS VDD net58 core.osr.next_result_w\[12\] net70 core.osr.result_r\[12\] VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_2123_ VSS VDD _1039_ _1410_ _0172_ VSS VDD sky130_fd_sc_hd__nor2_1
X_2054_ VSS VDD _1400_ _0133_ _1052_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_34_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_2956_ VSS VDD _0820_ _0848_ _0847_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1907_ VDD VSS _1377_ _1374_ _1376_ VSS VDD sky130_fd_sc_hd__and2_1
X_2887_ VSS VDD _0757_ _0781_ VSS VDD sky130_fd_sc_hd__clkbuf_2
X_1838_ VSS VDD _1326_ _1319_ _1327_ VSS VDD sky130_fd_sc_hd__nor2_1
X_1769_ VSS VDD _1249_ _1281_ _1213_ VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_103_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_103_146 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__2497__B1 _0439_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3120__RESET_B net85 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput52 VDD VSS result_out[8] net52 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput41 VDD VSS result_out[12] net41 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_48_200 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_56_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_2810_ VDD VSS _0705_ core.cnb.shift_register_r\[5\] VSS VDD sky130_fd_sc_hd__inv_2
X_2741_ VSS VDD net54 _0637_ core.cnb.is_holding_result_w VSS VDD sky130_fd_sc_hd__nor2_2
X_2672_ VSS VDD core.osr.next_result_w\[9\] _0575_ _0568_ VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1608__B _1045_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1623_ VDD VSS _1169_ _1128_ VSS VDD sky130_fd_sc_hd__inv_2
X_1554_ VSS VDD _1048_ _1108_ _1097_ VSS VDD sky130_fd_sc_hd__nand2_1
X_1485_ VSS VDD _1045_ core.cnb.data_register_r\[6\] core.cnb.data_register_r\[7\]
+ VSS VDD sky130_fd_sc_hd__nor2_4
.ends

.subckt adc_wrapper VDD rst_n clk conv_start conv_finish load dati dato tie0 tie1
+ inp_ana inn_ana VSS
Xadc_bridge_0 VDD adc_top_0/config_1_in[0] adc_top_0/config_1_in[10] adc_top_0/config_1_in[11]
+ adc_top_0/config_1_in[12] adc_top_0/config_1_in[13] adc_top_0/config_1_in[14] adc_top_0/config_1_in[15]
+ adc_top_0/config_1_in[1] adc_top_0/config_1_in[2] adc_top_0/config_1_in[3] adc_top_0/config_1_in[4]
+ adc_top_0/config_1_in[5] adc_top_0/config_1_in[6] adc_top_0/config_1_in[7] adc_top_0/config_1_in[8]
+ adc_top_0/config_1_in[9] adc_top_0/config_2_in[0] adc_top_0/config_2_in[10] adc_top_0/config_2_in[11]
+ adc_top_0/config_2_in[12] adc_top_0/config_2_in[13] adc_top_0/config_2_in[14] adc_top_0/config_2_in[15]
+ adc_top_0/config_2_in[1] adc_top_0/config_2_in[2] adc_top_0/config_2_in[3] adc_top_0/config_2_in[4]
+ adc_top_0/config_2_in[5] adc_top_0/config_2_in[6] adc_top_0/config_2_in[7] adc_top_0/config_2_in[8]
+ adc_top_0/config_2_in[9] adc_bridge_0/adc_conv_finished adc_bridge_0/adc_conv_finished_osr
+ adc_top_0/result_out[0] adc_top_0/result_out[10] adc_top_0/result_out[11] adc_top_0/result_out[12]
+ adc_top_0/result_out[13] adc_top_0/result_out[14] adc_top_0/result_out[15] adc_top_0/result_out[1]
+ adc_top_0/result_out[2] adc_top_0/result_out[3] adc_top_0/result_out[4] adc_top_0/result_out[5]
+ adc_top_0/result_out[6] adc_top_0/result_out[7] adc_top_0/result_out[8] adc_top_0/result_out[9]
+ clk conv_finish dati dato load rst_n tie0 tie1 VSS adc_bridge
Xadc_top_0 clk adc_top_0/config_1_in[0] adc_top_0/config_1_in[10] adc_top_0/config_1_in[11]
+ adc_top_0/config_1_in[12] adc_top_0/config_1_in[13] adc_top_0/config_1_in[14] adc_top_0/config_1_in[15]
+ adc_top_0/config_1_in[1] adc_top_0/config_1_in[2] adc_top_0/config_1_in[3] adc_top_0/config_1_in[4]
+ adc_top_0/config_1_in[5] adc_top_0/config_1_in[6] adc_top_0/config_1_in[7] adc_top_0/config_1_in[8]
+ adc_top_0/config_1_in[9] adc_top_0/config_2_in[0] adc_top_0/config_2_in[10] adc_top_0/config_2_in[11]
+ adc_top_0/config_2_in[12] adc_top_0/config_2_in[13] adc_top_0/config_2_in[14] adc_top_0/config_2_in[15]
+ adc_top_0/config_2_in[1] adc_top_0/config_2_in[2] adc_top_0/config_2_in[3] adc_top_0/config_2_in[4]
+ adc_top_0/config_2_in[5] adc_top_0/config_2_in[6] adc_top_0/config_2_in[7] adc_top_0/config_2_in[8]
+ adc_top_0/config_2_in[9] adc_bridge_0/adc_conv_finished_osr adc_bridge_0/adc_conv_finished
+ inn_ana inp_ana adc_top_0/result_out[0] adc_top_0/result_out[10] adc_top_0/result_out[11]
+ adc_top_0/result_out[12] adc_top_0/result_out[13] adc_top_0/result_out[14] adc_top_0/result_out[15]
+ adc_top_0/result_out[1] adc_top_0/result_out[2] adc_top_0/result_out[3] adc_top_0/result_out[4]
+ adc_top_0/result_out[5] adc_top_0/result_out[6] adc_top_0/result_out[7] adc_top_0/result_out[8]
+ adc_top_0/result_out[9] rst_n conv_start VDD VSS adc_top
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i io_analog[4]_uq0 io_analog[4]_uq1 io_analog[4]_uq2 io_analog[4]_uq3
+ io_analog[4]_uq4 io_analog[5]_uq0 io_analog[5]_uq1 io_analog[5]_uq2 io_analog[5]_uq3
+ io_analog[5]_uq4 io_analog[6]_uq0 io_analog[6]_uq1 io_analog[6]_uq2 io_analog[6]_uq3
+ io_analog[6]_uq4 vssa1_uq0 vssa1_uq1 vssa1_uq2 vssd2_uq0 vssa2_uq0 vdda2_uq0 vdda1_uq0
+ vdda1_uq1 vdda1_uq2 vccd2_uq0
Xmerg1b_0 io_analog[7] io_in[18] vdda2_uq0 io_analog[10] vssa2_uq0 io_analog[9] user_clock2
+ io_analog[8] io_in[19] io_in[25] io_in[20] io_out[24] io_in[17] merg1b
Xadc_wrapper_0 vccd1 io_in[11] io_in[13] io_in[12] io_out[5] io_in[8] io_in[7] io_out[6]
+ adc_wrapper_0/tie0 adc_wrapper_0/tie1 gpio_analog[3] gpio_analog[2] vssa2_uq0 adc_wrapper
R0 adc_wrapper_0/tie1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R1 adc_wrapper_0/tie1 io_oeb[13] sky130_fd_pr__res_generic_m3 w=0.3 l=0.59
R2 adc_wrapper_0/tie0 io_oeb[6] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R3 adc_wrapper_0/tie1 io_oeb[11] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R4 adc_wrapper_0/tie1 io_oeb[7] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R5 adc_wrapper_0/tie0 io_oeb[5] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R6 adc_wrapper_0/tie1 io_oeb[9] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R7 adc_wrapper_0/tie1 io_oeb[8] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
R8 adc_wrapper_0/tie1 io_oeb[10] sky130_fd_pr__res_generic_m3 w=0.3 l=0.6
.ends

