magic
tech sky130A
magscale 1 2
timestamp 1697806833
<< nwell >>
rect -3254 -3219 3254 3219
<< pmos >>
rect -3058 -3000 -1058 3000
rect -1000 -3000 1000 3000
rect 1058 -3000 3058 3000
<< pdiff >>
rect -3116 2988 -3058 3000
rect -3116 -2988 -3104 2988
rect -3070 -2988 -3058 2988
rect -3116 -3000 -3058 -2988
rect -1058 2988 -1000 3000
rect -1058 -2988 -1046 2988
rect -1012 -2988 -1000 2988
rect -1058 -3000 -1000 -2988
rect 1000 2988 1058 3000
rect 1000 -2988 1012 2988
rect 1046 -2988 1058 2988
rect 1000 -3000 1058 -2988
rect 3058 2988 3116 3000
rect 3058 -2988 3070 2988
rect 3104 -2988 3116 2988
rect 3058 -3000 3116 -2988
<< pdiffc >>
rect -3104 -2988 -3070 2988
rect -1046 -2988 -1012 2988
rect 1012 -2988 1046 2988
rect 3070 -2988 3104 2988
<< nsubdiff >>
rect -3218 3149 -3122 3183
rect 3122 3149 3218 3183
rect -3218 3087 -3184 3149
rect 3184 3087 3218 3149
rect -3218 -3149 -3184 -3087
rect 3184 -3149 3218 -3087
rect -3218 -3183 -3122 -3149
rect 3122 -3183 3218 -3149
<< nsubdiffcont >>
rect -3122 3149 3122 3183
rect -3218 -3087 -3184 3087
rect 3184 -3087 3218 3087
rect -3122 -3183 3122 -3149
<< poly >>
rect -3058 3081 -1058 3097
rect -3058 3047 -3042 3081
rect -1074 3047 -1058 3081
rect -3058 3000 -1058 3047
rect -1000 3081 1000 3097
rect -1000 3047 -984 3081
rect 984 3047 1000 3081
rect -1000 3000 1000 3047
rect 1058 3081 3058 3097
rect 1058 3047 1074 3081
rect 3042 3047 3058 3081
rect 1058 3000 3058 3047
rect -3058 -3047 -1058 -3000
rect -3058 -3081 -3042 -3047
rect -1074 -3081 -1058 -3047
rect -3058 -3097 -1058 -3081
rect -1000 -3047 1000 -3000
rect -1000 -3081 -984 -3047
rect 984 -3081 1000 -3047
rect -1000 -3097 1000 -3081
rect 1058 -3047 3058 -3000
rect 1058 -3081 1074 -3047
rect 3042 -3081 3058 -3047
rect 1058 -3097 3058 -3081
<< polycont >>
rect -3042 3047 -1074 3081
rect -984 3047 984 3081
rect 1074 3047 3042 3081
rect -3042 -3081 -1074 -3047
rect -984 -3081 984 -3047
rect 1074 -3081 3042 -3047
<< locali >>
rect -3218 3149 -3122 3183
rect 3122 3149 3218 3183
rect -3218 3087 -3184 3149
rect 3184 3087 3218 3149
rect -3058 3047 -3042 3081
rect -1074 3047 -1058 3081
rect -1000 3047 -984 3081
rect 984 3047 1000 3081
rect 1058 3047 1074 3081
rect 3042 3047 3058 3081
rect -3104 2988 -3070 3004
rect -3104 -3004 -3070 -2988
rect -1046 2988 -1012 3004
rect -1046 -3004 -1012 -2988
rect 1012 2988 1046 3004
rect 1012 -3004 1046 -2988
rect 3070 2988 3104 3004
rect 3070 -3004 3104 -2988
rect -3058 -3081 -3042 -3047
rect -1074 -3081 -1058 -3047
rect -1000 -3081 -984 -3047
rect 984 -3081 1000 -3047
rect 1058 -3081 1074 -3047
rect 3042 -3081 3058 -3047
rect -3218 -3149 -3184 -3087
rect 3184 -3149 3218 -3087
rect -3218 -3183 -3122 -3149
rect 3122 -3183 3218 -3149
<< viali >>
rect -3042 3047 -1074 3081
rect -984 3047 984 3081
rect 1074 3047 3042 3081
rect -3104 -2988 -3070 2988
rect -1046 -2988 -1012 2988
rect 1012 -2988 1046 2988
rect 3070 -2988 3104 2988
rect -3042 -3081 -1074 -3047
rect -984 -3081 984 -3047
rect 1074 -3081 3042 -3047
<< metal1 >>
rect -3054 3081 -1062 3087
rect -3054 3047 -3042 3081
rect -1074 3047 -1062 3081
rect -3054 3041 -1062 3047
rect -996 3081 996 3087
rect -996 3047 -984 3081
rect 984 3047 996 3081
rect -996 3041 996 3047
rect 1062 3081 3054 3087
rect 1062 3047 1074 3081
rect 3042 3047 3054 3081
rect 1062 3041 3054 3047
rect -3110 2988 -3064 3000
rect -3110 -2988 -3104 2988
rect -3070 -2988 -3064 2988
rect -3110 -3000 -3064 -2988
rect -1052 2988 -1006 3000
rect -1052 -2988 -1046 2988
rect -1012 -2988 -1006 2988
rect -1052 -3000 -1006 -2988
rect 1006 2988 1052 3000
rect 1006 -2988 1012 2988
rect 1046 -2988 1052 2988
rect 1006 -3000 1052 -2988
rect 3064 2988 3110 3000
rect 3064 -2988 3070 2988
rect 3104 -2988 3110 2988
rect 3064 -3000 3110 -2988
rect -3054 -3047 -1062 -3041
rect -3054 -3081 -3042 -3047
rect -1074 -3081 -1062 -3047
rect -3054 -3087 -1062 -3081
rect -996 -3047 996 -3041
rect -996 -3081 -984 -3047
rect 984 -3081 996 -3047
rect -996 -3087 996 -3081
rect 1062 -3047 3054 -3041
rect 1062 -3081 1074 -3047
rect 3042 -3081 3054 -3047
rect 1062 -3087 3054 -3081
<< properties >>
string FIXED_BBOX -3201 -3166 3201 3166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 30 l 10 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
