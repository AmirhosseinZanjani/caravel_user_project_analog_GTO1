magic
tech sky130A
magscale 1 2
timestamp 1698131850
use osc_nfet_w30_nf4_cc  osc_nfet_w30_nf4_cc_0
timestamp 1698131850
transform 1 0 10348 0 1 0
box 0 -240 5176 1957
use osc_nfet_w30_nf4_cc  osc_nfet_w30_nf4_cc_1
timestamp 1698131850
transform 1 0 5172 0 1 0
box 0 -240 5176 1957
<< end >>
