magic
tech sky130A
magscale 1 2
timestamp 1695810207
<< locali >>
rect -61 170 115 1170
rect 1589 170 1765 1170
rect 46 -4 86 132
rect 1618 -4 1658 132
<< metal1 >>
rect 204 1580 252 1584
rect 202 1574 254 1580
rect 202 1516 254 1522
rect 204 1170 252 1516
rect 300 1484 348 1584
rect 396 1580 444 1584
rect 394 1574 446 1580
rect 394 1516 446 1522
rect 298 1478 350 1484
rect 298 1420 350 1426
rect 300 1170 348 1420
rect 396 1170 444 1516
rect 492 1484 540 1584
rect 588 1580 636 1584
rect 586 1574 638 1580
rect 586 1516 638 1522
rect 490 1478 542 1484
rect 490 1420 542 1426
rect 492 1170 540 1420
rect 588 1170 636 1516
rect 684 1484 732 1584
rect 780 1580 828 1584
rect 778 1574 830 1580
rect 778 1516 830 1522
rect 682 1478 734 1484
rect 682 1420 734 1426
rect 684 1170 732 1420
rect 780 1170 828 1516
rect 876 1484 924 1584
rect 972 1580 1020 1584
rect 970 1574 1022 1580
rect 970 1516 1022 1522
rect 874 1478 926 1484
rect 874 1420 926 1426
rect 876 1170 924 1420
rect 972 1170 1020 1516
rect 1068 1484 1116 1584
rect 1164 1580 1212 1584
rect 1162 1574 1214 1580
rect 1162 1516 1214 1522
rect 1066 1478 1118 1484
rect 1066 1420 1118 1426
rect 1068 1170 1116 1420
rect 1164 1170 1212 1516
rect 1260 1484 1308 1584
rect 1356 1580 1404 1584
rect 1354 1574 1406 1580
rect 1354 1516 1406 1522
rect 1258 1478 1310 1484
rect 1258 1420 1310 1426
rect 1260 1170 1308 1420
rect 1356 1170 1404 1516
rect 1452 1484 1500 1584
rect 1450 1478 1502 1484
rect 1450 1420 1502 1426
rect 1452 1170 1500 1420
rect -131 91 1835 139
<< via1 >>
rect 202 1522 254 1574
rect 394 1522 446 1574
rect 298 1426 350 1478
rect 586 1522 638 1574
rect 490 1426 542 1478
rect 778 1522 830 1574
rect 682 1426 734 1478
rect 970 1522 1022 1574
rect 874 1426 926 1478
rect 1162 1522 1214 1574
rect 1066 1426 1118 1478
rect 1354 1522 1406 1574
rect 1258 1426 1310 1478
rect 1450 1426 1502 1478
<< metal2 >>
rect 202 1574 254 1580
rect -130 1524 202 1572
rect 394 1574 446 1580
rect 254 1524 394 1572
rect 202 1516 254 1522
rect 586 1574 638 1580
rect 446 1524 586 1572
rect 394 1516 446 1522
rect 778 1574 830 1580
rect 638 1524 778 1572
rect 586 1516 638 1522
rect 970 1574 1022 1580
rect 830 1524 970 1572
rect 778 1516 830 1522
rect 1162 1574 1214 1580
rect 1022 1524 1162 1572
rect 970 1516 1022 1522
rect 1354 1574 1406 1580
rect 1214 1524 1354 1572
rect 1162 1516 1214 1522
rect 1406 1524 1842 1572
rect 1354 1516 1406 1522
rect 298 1478 350 1484
rect -130 1428 298 1476
rect 490 1478 542 1484
rect 350 1428 490 1476
rect 298 1420 350 1426
rect 682 1478 734 1484
rect 542 1428 682 1476
rect 490 1420 542 1426
rect 874 1478 926 1484
rect 734 1428 874 1476
rect 682 1420 734 1426
rect 1066 1478 1118 1484
rect 926 1428 1066 1476
rect 874 1420 926 1426
rect 1258 1478 1310 1484
rect 1118 1428 1258 1476
rect 1066 1420 1118 1426
rect 1450 1478 1502 1484
rect 1310 1428 1450 1476
rect 1258 1420 1310 1426
rect 1502 1428 1842 1476
rect 1450 1420 1502 1426
use sky130_fd_pr__nfet_01v8_YN9FL4  sky130_fd_pr__nfet_01v8_UDPJLN_0
timestamp 1695643842
transform 1 0 852 0 1 670
box -983 -710 983 710
<< labels >>
flabel locali -61 170 115 1170 0 FreeSans 240 0 0 0 vss_sw
port 0 nsew
flabel metal2 -130 1524 202 1572 0 FreeSans 240 0 0 0 vp_sw
port 2 nsew
flabel metal2 -130 1428 202 1476 0 FreeSans 240 0 0 0 vn_sw
port 3 nsew
flabel metal1 -131 91 1835 139 0 FreeSans 240 0 0 0 en_sw
port 1 nsew
<< end >>
