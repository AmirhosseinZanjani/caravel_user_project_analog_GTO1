magic
tech sky130A
magscale 1 2
timestamp 1698131850
<< locali >>
rect 3761 25870 4079 26006
rect 6749 25870 7067 26006
rect 3667 25082 4173 25832
rect 6655 25082 7161 25832
rect 11947 24243 17512 25910
rect 22428 25870 22746 26006
rect 25416 25870 25734 26006
rect 22334 25082 22840 25832
rect 25322 25082 25828 25832
rect 11947 22090 17512 22963
rect 14559 21329 14763 22090
<< metal1 >>
rect 2826 27396 2878 27402
rect 2826 27194 2878 27200
rect 3162 27396 3214 27402
rect 3162 27194 3214 27200
rect 26281 27396 26333 27402
rect 26281 27194 26333 27200
rect 26617 27396 26669 27402
rect 26617 27194 26669 27200
rect 2828 26188 2876 27194
rect 3164 26188 3212 27194
rect 4628 27106 4676 27122
rect 4964 27106 5012 27122
rect 5816 27106 5864 27122
rect 6152 27106 6200 27122
rect 23295 27106 23343 27122
rect 23631 27106 23679 27122
rect 24483 27106 24531 27122
rect 24819 27106 24867 27122
rect 4626 27100 4678 27106
rect 4626 26898 4678 26904
rect 4962 27100 5014 27106
rect 4962 26898 5014 26904
rect 5814 27100 5866 27106
rect 5814 26898 5866 26904
rect 6150 27100 6202 27106
rect 6150 26898 6202 26904
rect 23294 27100 23346 27106
rect 23294 26898 23346 26904
rect 23630 27100 23682 27106
rect 23630 26898 23682 26904
rect 24482 27100 24534 27106
rect 24482 26898 24534 26904
rect 24818 27100 24870 27106
rect 24818 26898 24870 26904
rect 4628 26188 4676 26898
rect 4964 26188 5012 26898
rect 5816 26233 5864 26898
rect 6152 26188 6200 26898
rect 23295 26188 23343 26898
rect 23631 26233 23679 26898
rect 24483 26194 24531 26898
rect 24819 26188 24867 26898
rect 26283 26188 26331 27194
rect 26619 26188 26667 27194
rect -6712 -16158 15550 -16128
rect -6712 -16698 -6681 -16158
rect -3931 -16698 15550 -16158
rect -6712 -17128 15550 -16698
rect -6711 -21830 15550 -21400
rect -6711 -22370 -6681 -21830
rect -3931 -22370 15550 -21830
rect -6711 -22400 15550 -22370
rect 13950 -27982 15550 -24905
rect -6712 -28012 15550 -27982
rect -6712 -28552 -6681 -28012
rect -3931 -28552 15550 -28012
rect -6712 -28982 15550 -28552
rect 13950 -33254 15550 -28982
rect -6711 -33684 15550 -33254
rect -6711 -34224 -6681 -33684
rect -3931 -34224 15550 -33684
rect -6711 -34254 15550 -34224
<< via1 >>
rect 2826 27200 2878 27396
rect 3162 27200 3214 27396
rect 26281 27200 26333 27396
rect 26617 27200 26669 27396
rect 4626 26904 4678 27100
rect 4962 26904 5014 27100
rect 5814 26904 5866 27100
rect 6150 26904 6202 27100
rect 23294 26904 23346 27100
rect 23630 26904 23682 27100
rect 24482 26904 24534 27100
rect 24818 26904 24870 27100
rect -6681 -16698 -3931 -16158
rect -6681 -22370 -3931 -21830
rect -6681 -28552 -3931 -28012
rect -6681 -34224 -3931 -33684
<< metal2 >>
rect 2826 27396 2878 27402
rect 2373 27202 2826 27394
rect 3162 27396 3214 27402
rect 2878 27202 3162 27394
rect 2826 27194 2878 27200
rect 26281 27396 26333 27402
rect 3214 27202 26281 27394
rect 3162 27194 3214 27200
rect 26617 27396 26669 27402
rect 26333 27202 26617 27394
rect 26281 27194 26333 27200
rect 26669 27202 27122 27394
rect 26617 27194 26669 27200
rect 4626 27100 4678 27106
rect 2373 26906 4626 27098
rect 4962 27100 5014 27106
rect 4678 26906 4962 27098
rect 4626 26898 4678 26904
rect 5814 27100 5866 27106
rect 5014 26906 5814 27098
rect 4962 26898 5014 26904
rect 6150 27100 6202 27106
rect 5866 26906 6150 27098
rect 5814 26898 5866 26904
rect 23294 27100 23346 27106
rect 6202 26906 23294 27098
rect 6150 26898 6202 26904
rect 23630 27100 23682 27106
rect 23346 26906 23630 27098
rect 23294 26898 23346 26904
rect 24482 27100 24534 27106
rect 23682 26906 24482 27098
rect 23630 26898 23682 26904
rect 24818 27100 24870 27106
rect 24534 26906 24818 27098
rect 24482 26898 24534 26904
rect 24870 26906 27122 27098
rect 24818 26898 24870 26904
rect 2373 26744 12019 26804
rect 2373 26294 2433 26744
rect 7159 26294 12019 26744
rect 2373 26234 12019 26294
rect 17476 26745 27122 26804
rect 17476 26294 22335 26745
rect 27062 26294 27122 26745
rect 17476 26234 27122 26294
rect 7161 25994 22412 26186
rect 25322 26090 25407 26186
rect 27122 26090 27207 26186
rect 2373 24476 12019 24536
rect 2373 24026 2433 24476
rect 10903 24026 12019 24476
rect 2373 23966 12019 24026
rect 17476 24476 27122 24536
rect 17476 24026 18592 24476
rect 26989 24026 27122 24476
rect 17476 23966 27122 24026
rect 2373 23752 11983 23812
rect 2373 23302 2433 23752
rect 7159 23302 11983 23752
rect 2373 23242 11983 23302
rect 17512 23752 27122 23812
rect 17512 23302 22335 23752
rect 27062 23302 27122 23752
rect 17512 23242 27122 23302
rect 2373 23002 27198 23194
rect 2373 21484 11288 21544
rect 17512 21484 27122 21544
rect 2373 21034 2433 21484
rect 10867 21456 11959 21484
rect 10867 21034 11983 21456
rect 2373 20974 11983 21034
rect 17512 21034 18628 21484
rect 27062 21034 27122 21484
rect 17512 20974 27122 21034
rect -6712 -16158 -3902 -16128
rect -6712 -16698 -6681 -16158
rect -3931 -16698 -3902 -16158
rect -6712 -17128 -3902 -16698
rect -6711 -21830 -3901 -21400
rect -6711 -22370 -6681 -21830
rect -3931 -22370 -3901 -21830
rect -6711 -22400 -3901 -22370
rect -6712 -28012 -3902 -27982
rect -6712 -28552 -6681 -28012
rect -3931 -28552 -3902 -28012
rect -6712 -28982 -3902 -28552
rect -6711 -33684 -3901 -33254
rect -6711 -34224 -6681 -33684
rect -3931 -34224 -3901 -33684
rect -6711 -34254 -3901 -34224
<< via2 >>
rect 2433 26294 7159 26744
rect 22335 26294 27062 26745
rect 2433 24026 10903 24476
rect 18592 24026 26989 24476
rect 2433 23302 7159 23752
rect 22335 23302 27062 23752
rect 2433 21034 10867 21484
rect 18628 21034 27062 21484
rect -6681 -16698 -3931 -16158
rect -6681 -22370 -3931 -21830
rect -6681 -28552 -3931 -28012
rect -6681 -34224 -3931 -33684
<< metal3 >>
rect 2373 26744 7219 26804
rect 2373 26294 2433 26744
rect 7159 26294 7219 26744
rect 2373 26234 7219 26294
rect 22275 26745 27122 26804
rect 22275 26294 22335 26745
rect 27062 26294 27122 26745
rect 22275 26234 27122 26294
rect 2373 24476 12019 24536
rect 2373 24026 2433 24476
rect 10903 24026 12019 24476
rect 2373 23966 12019 24026
rect 17476 24476 27122 24536
rect 17476 24026 18592 24476
rect 27062 24026 27122 24476
rect 17476 23966 27122 24026
rect 2373 23752 7219 23812
rect 2373 23302 2433 23752
rect 7159 23302 7219 23752
rect 2373 23242 7219 23302
rect 22275 23752 27122 23812
rect 22275 23302 22335 23752
rect 27062 23302 27122 23752
rect 22275 23242 27122 23302
rect 2373 21484 11288 21544
rect 17476 21484 27122 21544
rect 2373 21034 2433 21484
rect 10867 21456 11959 21484
rect 10867 21034 11983 21456
rect 2373 20974 11983 21034
rect 17476 21034 18628 21484
rect 27062 21034 27122 21484
rect 17476 20974 27122 21034
rect -6712 -16158 -3902 -16128
rect -6712 -16698 -6681 -16158
rect -3931 -16698 -3902 -16158
rect -6712 -16728 -3902 -16698
rect -6711 -21830 -3901 -21800
rect -6711 -22370 -6681 -21830
rect -3931 -22370 -3901 -21830
rect -6711 -22400 -3901 -22370
rect -6712 -28012 -3902 -27982
rect -6712 -28552 -6681 -28012
rect -3931 -28552 -3902 -28012
rect -6712 -28582 -3902 -28552
rect -6711 -33684 -3901 -33654
rect -6711 -34224 -6681 -33684
rect -3931 -34224 -3901 -33684
rect -6711 -34254 -3901 -34224
<< via3 >>
rect 2433 26294 7159 26744
rect 22335 26294 27062 26745
rect 2433 24026 10903 24476
rect 18592 24026 26989 24476
rect 26989 24026 27062 24476
rect 2433 23302 7159 23752
rect 22335 23302 27062 23752
rect 2433 21034 10867 21484
rect 18628 21034 27062 21484
rect -6681 -16698 -3931 -16158
rect -6681 -22370 -3931 -21830
rect -6681 -28552 -3931 -28012
rect -6681 -34224 -3931 -33684
<< metal4 >>
rect 2372 29446 27122 29506
rect 2372 28996 17535 29446
rect 18416 28996 23836 29446
rect 24716 28996 27122 29446
rect 2372 28936 27122 28996
rect 2373 28748 27122 28808
rect 2373 28298 4778 28748
rect 5658 28298 11079 28748
rect 11960 28298 27122 28748
rect 2373 28238 27122 28298
rect 8044 27468 21450 27528
rect 8044 27018 17534 27468
rect 18415 27018 21450 27468
rect 8044 26958 21450 27018
rect 2373 26744 7219 26804
rect 2373 26294 2433 26744
rect 7159 26294 7219 26744
rect 2373 26234 7219 26294
rect 22275 26745 27122 26804
rect 22275 26294 22335 26745
rect 27062 26294 27122 26745
rect 22275 26234 27122 26294
rect 8044 25846 21450 25906
rect 8044 25396 11079 25846
rect 11960 25396 21450 25846
rect 8044 25336 21450 25396
rect 2373 24476 12019 24536
rect 2373 24026 2433 24476
rect 10903 24026 12019 24476
rect 2373 23966 12019 24026
rect 17476 24476 27122 24536
rect 17476 24026 18592 24476
rect 27062 24026 27122 24476
rect 17476 23966 27122 24026
rect 2373 23752 7219 23812
rect 2373 23302 2433 23752
rect 7159 23302 7219 23752
rect 2373 23242 7219 23302
rect 22275 23752 27122 23812
rect 22275 23302 22335 23752
rect 27062 23302 27122 23752
rect 22275 23242 27122 23302
rect 2373 21484 12019 21544
rect 2373 21034 2433 21484
rect 10867 21034 12019 21484
rect 2373 20974 12019 21034
rect 17476 21484 27122 21544
rect 17476 21034 18628 21484
rect 27062 21034 27122 21484
rect 17476 20974 27122 21034
rect -6712 -16158 -3902 -16128
rect -6712 -16698 -6681 -16158
rect -3931 -16698 -3902 -16158
rect -6712 -17128 -3902 -16698
rect -6711 -19029 -3901 -18779
rect -6711 -19528 -6621 -19029
rect -3991 -19528 -3901 -19029
rect -6711 -19779 -3901 -19528
rect -6711 -21830 -3901 -21400
rect -6711 -22370 -6681 -21830
rect -3931 -22370 -3901 -21830
rect -6711 -22400 -3901 -22370
rect -6712 -28012 -3902 -27982
rect -6712 -28552 -6681 -28012
rect -3931 -28552 -3902 -28012
rect -6712 -28982 -3902 -28552
rect -6711 -30883 -3901 -30633
rect -6711 -31382 -6621 -30883
rect -3991 -31382 -3901 -30883
rect -6711 -31633 -3901 -31382
rect -6711 -33684 -3901 -33254
rect -6711 -34224 -6681 -33684
rect -3931 -34224 -3901 -33684
rect -6711 -34254 -3901 -34224
<< via4 >>
rect 17535 28996 18416 29446
rect 23836 28996 24716 29446
rect 4778 28298 5658 28748
rect 11079 28298 11960 28748
rect 17534 27018 18415 27468
rect 4778 26294 5658 26744
rect 23836 26294 24716 26744
rect 11079 25396 11960 25846
rect 4778 23302 5658 23752
rect 23836 23302 24716 23752
rect -6621 -19528 -3991 -19029
rect -6621 -31382 -3991 -30883
<< metal5 >>
rect 4718 28748 5718 29506
rect 4718 28298 4778 28748
rect 5658 28298 5718 28748
rect 4718 26744 5718 28298
rect 11019 28748 12019 32036
rect 11019 28298 11079 28748
rect 11960 28298 12019 28748
rect 11019 28238 12019 28298
rect 17475 29446 18475 32036
rect 17475 28996 17535 29446
rect 18416 28996 18475 29446
rect 17475 28238 18475 28996
rect 23776 29446 24776 29506
rect 23776 28996 23836 29446
rect 24716 28996 24776 29446
rect 4718 26294 4778 26744
rect 5658 26294 5718 26744
rect 4718 23752 5718 26294
rect 4718 23302 4778 23752
rect 5658 23302 5718 23752
rect 4718 23242 5718 23302
rect 11019 25846 12019 27661
rect 11019 25396 11079 25846
rect 11960 25396 12019 25846
rect 11019 -7940 12019 25396
rect 17475 27468 18475 27663
rect 17475 27018 17534 27468
rect 18415 27018 18475 27468
rect 17475 -7940 18475 27018
rect 23776 26744 24776 28996
rect 23776 26294 23836 26744
rect 24716 26294 24776 26744
rect 23776 23752 24776 26294
rect 23776 23302 23836 23752
rect 24716 23302 24776 23752
rect 23776 23242 24776 23302
rect 14247 -8504 15247 -8312
rect -8711 -19029 -3267 -18779
rect -8711 -19528 -6621 -19029
rect -3991 -19528 -3267 -19029
rect -8711 -19779 -3267 -19528
rect -8711 -30883 -3267 -30633
rect -8711 -31382 -6621 -30883
rect -3991 -31382 -3267 -30883
rect -8711 -31633 -3267 -31382
use balun  balun_0
timestamp 1698088655
transform 0 1 -37253 1 0 -25206
box -16698 33886 17366 69252
use pa_nfet_w15_nf4  pa_nfet_w15_nf4_0
timestamp 1697705955
transform -1 0 26988 0 -1 26020
box -134 -318 1160 1588
use pa_nfet_w15_nf4  pa_nfet_w15_nf4_1
timestamp 1697705955
transform 1 0 2507 0 -1 26020
box -134 -318 1160 1588
use pa_nfet_w30_nf4  pa_nfet_w30_nf4_0
timestamp 1698131850
transform 1 0 4227 0 -1 26253
box -54 -85 2428 1821
use pa_nfet_w30_nf4  pa_nfet_w30_nf4_1
timestamp 1698131850
transform -1 0 25268 0 -1 26253
box -54 -85 2428 1821
use pa_nfet_w60_nf4  pa_nfet_w60_nf4_0
timestamp 1698131850
transform -1 0 22334 0 -1 26245
box 0 -93 4858 1813
use pa_nfet_w60_nf4  pa_nfet_w60_nf4_2
timestamp 1698131850
transform 1 0 7161 0 -1 26245
box 0 -93 4858 1813
use pa_nfet_w120_nf4  pa_nfet_w120_nf4_0
timestamp 1698131850
transform 1 0 17512 0 -1 23253
box 0 -93 9610 1813
use pa_nfet_w120_nf4  pa_nfet_w120_nf4_1
timestamp 1698131850
transform 1 0 2373 0 -1 23253
box 0 -93 9610 1813
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_64
timestamp 1696250317
transform 0 1 18000 1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_65
timestamp 1696250317
transform 0 1 16570 -1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_70
timestamp 1696250317
transform 0 -1 11494 -1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_71
timestamp 1696250317
transform 0 1 12924 1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_0
timestamp 1698080665
transform 0 -1 -6071 -1 0 -32458
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_1
timestamp 1698080665
transform 0 -1 -4541 1 0 -32458
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_2
timestamp 1698080665
transform 0 -1 -4541 -1 0 -29807
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_3
timestamp 1698080665
transform 0 -1 -6071 1 0 -29807
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_4
timestamp 1698080665
transform 0 -1 -6071 -1 0 -20604
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_5
timestamp 1698080665
transform 0 -1 -4541 1 0 -20604
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_6
timestamp 1698080665
transform 0 -1 -4541 -1 0 -17953
box -986 -640 986 640
use sky130_fd_pr__cap_mim_m3_1_WE7GNF  sky130_fd_pr__cap_mim_m3_1_WE7GNF_7
timestamp 1698080665
transform 0 -1 -6071 1 0 -17953
box -986 -640 986 640
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_0
timestamp 1696579262
transform 1 0 3920 0 -1 25457
box -359 -585 359 585
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_1
timestamp 1696579262
transform 1 0 6908 0 -1 25457
box -359 -585 359 585
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_2
timestamp 1696579262
transform -1 0 22587 0 -1 25457
box -359 -585 359 585
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_3
timestamp 1696579262
transform -1 0 25575 0 -1 25457
box -359 -585 359 585
<< labels >>
flabel locali 14559 21329 14763 22090 0 FreeSans 1600 0 0 0 vss_pa
port 0 nsew
flabel metal2 27122 23098 27198 23194 0 FreeSans 320 0 0 0 en_pa[3]
port 3 nsew
flabel metal2 22334 26090 22412 26186 0 FreeSans 320 0 0 0 en_pa[2]
port 4 nsew
flabel metal2 25322 26090 25407 26186 0 FreeSans 320 0 0 0 en_pa[1]
port 5 nsew
flabel metal2 27122 26090 27207 26186 0 FreeSans 320 0 0 0 en_pa[0]
port 6 nsew
flabel metal5 17475 -7940 18475 -7176 0 FreeSans 1600 0 0 0 tunep_pa
port 7 nsew
flabel metal5 11019 -7940 12019 -7176 0 FreeSans 1600 0 0 0 tunen_pa
port 8 nsew
flabel metal5 11019 28748 12019 32036 0 FreeSans 1600 0 0 0 inn_pa
port 2 nsew
flabel metal5 17475 29446 18475 32036 0 FreeSans 1600 0 0 0 inp_pa
port 1 nsew
flabel metal5 -8711 -19779 -6621 -18779 0 FreeSans 1600 0 0 0 outp_pa
port 9 nsew
flabel metal5 -8711 -31633 -6621 -30633 0 FreeSans 1600 0 0 0 outn_pa
port 10 nsew
flabel metal5 14247 -8504 15247 -8312 0 FreeSans 1600 0 0 0 vdd_pa
port 11 nsew
<< end >>
