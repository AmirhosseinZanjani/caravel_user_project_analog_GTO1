magic
tech sky130A
magscale 1 2
timestamp 1699608013
<< viali >>
rect 2697 77469 2731 77503
rect 2881 77401 2915 77435
rect 8217 74205 8251 74239
rect 8401 74069 8435 74103
rect 6377 73729 6411 73763
rect 6745 73661 6779 73695
rect 7021 73661 7055 73695
rect 6561 73525 6595 73559
rect 8493 73525 8527 73559
rect 7757 73321 7791 73355
rect 7113 73185 7147 73219
rect 5089 73117 5123 73151
rect 7297 73117 7331 73151
rect 7941 73117 7975 73151
rect 5365 73049 5399 73083
rect 8125 73049 8159 73083
rect 6837 72981 6871 73015
rect 7205 72981 7239 73015
rect 7665 72981 7699 73015
rect 8217 72981 8251 73015
rect 5457 72777 5491 72811
rect 6377 72777 6411 72811
rect 5641 72641 5675 72675
rect 6745 72641 6779 72675
rect 7389 72641 7423 72675
rect 6837 72573 6871 72607
rect 6929 72573 6963 72607
rect 7205 72437 7239 72471
rect 4813 72097 4847 72131
rect 6745 72097 6779 72131
rect 7021 72097 7055 72131
rect 5089 71961 5123 71995
rect 6561 71893 6595 71927
rect 8493 71893 8527 71927
rect 5273 71689 5307 71723
rect 6377 71689 6411 71723
rect 6745 71689 6779 71723
rect 7205 71689 7239 71723
rect 8401 71689 8435 71723
rect 7573 71621 7607 71655
rect 8125 71621 8159 71655
rect 5457 71553 5491 71587
rect 7665 71553 7699 71587
rect 6837 71485 6871 71519
rect 6929 71485 6963 71519
rect 7849 71485 7883 71519
rect 6101 71009 6135 71043
rect 5365 70941 5399 70975
rect 5917 70941 5951 70975
rect 7205 70941 7239 70975
rect 8217 70941 8251 70975
rect 5181 70805 5215 70839
rect 5549 70805 5583 70839
rect 6009 70805 6043 70839
rect 7021 70805 7055 70839
rect 8401 70805 8435 70839
rect 4721 70533 4755 70567
rect 7021 70533 7055 70567
rect 4445 70465 4479 70499
rect 6745 70465 6779 70499
rect 6193 70397 6227 70431
rect 8493 70397 8527 70431
rect 6929 70057 6963 70091
rect 7573 69921 7607 69955
rect 7297 69853 7331 69887
rect 7389 69717 7423 69751
rect 4445 69377 4479 69411
rect 7205 69377 7239 69411
rect 8217 69377 8251 69411
rect 4721 69309 4755 69343
rect 6193 69309 6227 69343
rect 7297 69309 7331 69343
rect 7481 69309 7515 69343
rect 6837 69173 6871 69207
rect 8401 69173 8435 69207
rect 5181 68969 5215 69003
rect 8493 68969 8527 69003
rect 6009 68833 6043 68867
rect 6193 68833 6227 68867
rect 5365 68765 5399 68799
rect 5917 68765 5951 68799
rect 6469 68765 6503 68799
rect 6745 68765 6779 68799
rect 7021 68697 7055 68731
rect 5549 68629 5583 68663
rect 6653 68629 6687 68663
rect 5457 68425 5491 68459
rect 5825 68425 5859 68459
rect 5365 68289 5399 68323
rect 5917 68289 5951 68323
rect 7113 68289 7147 68323
rect 7205 68289 7239 68323
rect 8217 68289 8251 68323
rect 6101 68221 6135 68255
rect 7021 68221 7055 68255
rect 5181 68085 5215 68119
rect 7573 68085 7607 68119
rect 8401 68085 8435 68119
rect 6561 67881 6595 67915
rect 8493 67881 8527 67915
rect 4813 67745 4847 67779
rect 5089 67745 5123 67779
rect 6745 67677 6779 67711
rect 7021 67609 7055 67643
rect 6745 67337 6779 67371
rect 7205 67337 7239 67371
rect 6837 67269 6871 67303
rect 7389 67201 7423 67235
rect 8217 67201 8251 67235
rect 6929 67133 6963 67167
rect 6377 66997 6411 67031
rect 8401 66997 8435 67031
rect 6561 66793 6595 66827
rect 4813 66657 4847 66691
rect 8125 66657 8159 66691
rect 8217 66657 8251 66691
rect 5089 66521 5123 66555
rect 6653 66521 6687 66555
rect 7389 66521 7423 66555
rect 8033 66521 8067 66555
rect 7665 66453 7699 66487
rect 5273 66249 5307 66283
rect 8493 66249 8527 66283
rect 5457 66113 5491 66147
rect 6469 66113 6503 66147
rect 6745 66045 6779 66079
rect 7021 66045 7055 66079
rect 6653 65977 6687 66011
rect 4813 65569 4847 65603
rect 7481 65569 7515 65603
rect 7297 65501 7331 65535
rect 8217 65501 8251 65535
rect 5089 65433 5123 65467
rect 6837 65433 6871 65467
rect 6929 65365 6963 65399
rect 7389 65365 7423 65399
rect 8401 65365 8435 65399
rect 5641 65161 5675 65195
rect 4721 65093 4755 65127
rect 8125 65093 8159 65127
rect 5549 65025 5583 65059
rect 5825 65025 5859 65059
rect 6837 65025 6871 65059
rect 7021 64821 7055 64855
rect 8217 64821 8251 64855
rect 7021 64481 7055 64515
rect 6469 64413 6503 64447
rect 6745 64413 6779 64447
rect 6653 64277 6687 64311
rect 8493 64277 8527 64311
rect 5273 64073 5307 64107
rect 6745 64005 6779 64039
rect 4997 63937 5031 63971
rect 5641 63937 5675 63971
rect 5733 63869 5767 63903
rect 5825 63869 5859 63903
rect 6469 63869 6503 63903
rect 4813 63733 4847 63767
rect 8217 63733 8251 63767
rect 4616 63529 4650 63563
rect 6101 63529 6135 63563
rect 6377 63529 6411 63563
rect 7205 63461 7239 63495
rect 8401 63461 8435 63495
rect 4353 63393 4387 63427
rect 6837 63393 6871 63427
rect 7021 63393 7055 63427
rect 7849 63393 7883 63427
rect 6745 63325 6779 63359
rect 8125 63325 8159 63359
rect 7573 63257 7607 63291
rect 7665 63189 7699 63223
rect 5549 62985 5583 63019
rect 4997 62849 5031 62883
rect 5641 62849 5675 62883
rect 8217 62849 8251 62883
rect 5825 62781 5859 62815
rect 5181 62713 5215 62747
rect 4813 62645 4847 62679
rect 8401 62645 8435 62679
rect 4353 62305 4387 62339
rect 4629 62305 4663 62339
rect 6469 62237 6503 62271
rect 6745 62237 6779 62271
rect 7021 62169 7055 62203
rect 6101 62101 6135 62135
rect 6653 62101 6687 62135
rect 8493 62101 8527 62135
rect 6745 61897 6779 61931
rect 7113 61897 7147 61931
rect 7205 61829 7239 61863
rect 7389 61693 7423 61727
rect 4445 61217 4479 61251
rect 6837 61149 6871 61183
rect 8217 61149 8251 61183
rect 4721 61081 4755 61115
rect 7481 61081 7515 61115
rect 6193 61013 6227 61047
rect 7021 61013 7055 61047
rect 7389 61013 7423 61047
rect 8401 61013 8435 61047
rect 4813 60809 4847 60843
rect 5549 60809 5583 60843
rect 7021 60741 7055 60775
rect 4997 60673 5031 60707
rect 5641 60673 5675 60707
rect 5825 60605 5859 60639
rect 6745 60605 6779 60639
rect 5181 60537 5215 60571
rect 8493 60469 8527 60503
rect 6653 60265 6687 60299
rect 5181 60197 5215 60231
rect 5825 60129 5859 60163
rect 7205 60129 7239 60163
rect 5089 60061 5123 60095
rect 7021 60061 7055 60095
rect 8217 60061 8251 60095
rect 5549 59993 5583 60027
rect 7113 59993 7147 60027
rect 4905 59925 4939 59959
rect 5641 59925 5675 59959
rect 8401 59925 8435 59959
rect 6653 59721 6687 59755
rect 4721 59653 4755 59687
rect 7021 59653 7055 59687
rect 4445 59585 4479 59619
rect 6469 59585 6503 59619
rect 6745 59517 6779 59551
rect 6193 59381 6227 59415
rect 8493 59381 8527 59415
rect 6745 59177 6779 59211
rect 5917 59041 5951 59075
rect 7205 59041 7239 59075
rect 7389 59041 7423 59075
rect 5641 58973 5675 59007
rect 7113 58973 7147 59007
rect 8125 58905 8159 58939
rect 5273 58837 5307 58871
rect 5733 58837 5767 58871
rect 8401 58837 8435 58871
rect 4721 58565 4755 58599
rect 6469 58497 6503 58531
rect 4445 58429 4479 58463
rect 6745 58429 6779 58463
rect 7021 58429 7055 58463
rect 6653 58361 6687 58395
rect 6193 58293 6227 58327
rect 8493 58293 8527 58327
rect 4997 58089 5031 58123
rect 6745 58089 6779 58123
rect 7389 57953 7423 57987
rect 5181 57885 5215 57919
rect 7113 57885 7147 57919
rect 8125 57817 8159 57851
rect 7205 57749 7239 57783
rect 8217 57749 8251 57783
rect 6837 57409 6871 57443
rect 7757 57409 7791 57443
rect 4445 57341 4479 57375
rect 4721 57341 4755 57375
rect 6193 57205 6227 57239
rect 7021 57205 7055 57239
rect 8033 57205 8067 57239
rect 4813 57001 4847 57035
rect 6009 57001 6043 57035
rect 5089 56933 5123 56967
rect 6377 56933 6411 56967
rect 5733 56865 5767 56899
rect 6745 56865 6779 56899
rect 7021 56865 7055 56899
rect 8493 56865 8527 56899
rect 4997 56797 5031 56831
rect 5457 56797 5491 56831
rect 6193 56797 6227 56831
rect 5549 56661 5583 56695
rect 5273 56457 5307 56491
rect 6561 56457 6595 56491
rect 6745 56457 6779 56491
rect 7113 56457 7147 56491
rect 5641 56389 5675 56423
rect 7205 56389 7239 56423
rect 5181 56321 5215 56355
rect 6469 56321 6503 56355
rect 5733 56253 5767 56287
rect 5917 56253 5951 56287
rect 7297 56253 7331 56287
rect 4997 56117 5031 56151
rect 4813 55777 4847 55811
rect 6745 55777 6779 55811
rect 4537 55709 4571 55743
rect 6469 55709 6503 55743
rect 7021 55641 7055 55675
rect 6285 55573 6319 55607
rect 6653 55573 6687 55607
rect 8493 55573 8527 55607
rect 6653 55369 6687 55403
rect 7113 55301 7147 55335
rect 7021 55233 7055 55267
rect 7849 55233 7883 55267
rect 8493 55233 8527 55267
rect 7205 55165 7239 55199
rect 7573 54825 7607 54859
rect 4537 54621 4571 54655
rect 8217 54621 8251 54655
rect 4813 54553 4847 54587
rect 7665 54553 7699 54587
rect 6285 54485 6319 54519
rect 8401 54485 8435 54519
rect 4997 54281 5031 54315
rect 5273 54281 5307 54315
rect 5641 54281 5675 54315
rect 5181 54145 5215 54179
rect 6469 54145 6503 54179
rect 6745 54145 6779 54179
rect 5733 54077 5767 54111
rect 5917 54077 5951 54111
rect 7021 54077 7055 54111
rect 6653 54009 6687 54043
rect 8493 53941 8527 53975
rect 6653 53737 6687 53771
rect 5917 53601 5951 53635
rect 7205 53601 7239 53635
rect 5181 53533 5215 53567
rect 7021 53533 7055 53567
rect 5641 53465 5675 53499
rect 7113 53465 7147 53499
rect 4997 53397 5031 53431
rect 5273 53397 5307 53431
rect 5733 53397 5767 53431
rect 4721 53125 4755 53159
rect 6469 53057 6503 53091
rect 6745 53057 6779 53091
rect 4445 52989 4479 53023
rect 7021 52989 7055 53023
rect 6653 52921 6687 52955
rect 6193 52853 6227 52887
rect 8493 52853 8527 52887
rect 6653 52649 6687 52683
rect 8401 52649 8435 52683
rect 7113 52513 7147 52547
rect 7205 52513 7239 52547
rect 7021 52445 7055 52479
rect 8217 52445 8251 52479
rect 8217 51969 8251 52003
rect 4445 51901 4479 51935
rect 4721 51901 4755 51935
rect 6193 51765 6227 51799
rect 8401 51765 8435 51799
rect 4905 51561 4939 51595
rect 5733 51425 5767 51459
rect 5917 51425 5951 51459
rect 6745 51425 6779 51459
rect 5089 51357 5123 51391
rect 5641 51357 5675 51391
rect 6469 51357 6503 51391
rect 7021 51289 7055 51323
rect 5273 51221 5307 51255
rect 6653 51221 6687 51255
rect 8493 51221 8527 51255
rect 5365 51017 5399 51051
rect 6653 51017 6687 51051
rect 7021 51017 7055 51051
rect 5181 50881 5215 50915
rect 5733 50881 5767 50915
rect 7113 50881 7147 50915
rect 5825 50813 5859 50847
rect 5917 50813 5951 50847
rect 7205 50813 7239 50847
rect 4997 50677 5031 50711
rect 6285 50473 6319 50507
rect 6653 50405 6687 50439
rect 4813 50337 4847 50371
rect 7021 50337 7055 50371
rect 4537 50269 4571 50303
rect 6469 50269 6503 50303
rect 6745 50269 6779 50303
rect 8493 50133 8527 50167
rect 8401 49929 8435 49963
rect 5457 49793 5491 49827
rect 7481 49793 7515 49827
rect 8217 49793 8251 49827
rect 4629 49725 4663 49759
rect 6653 49725 6687 49759
rect 6653 49385 6687 49419
rect 7205 49249 7239 49283
rect 4721 49181 4755 49215
rect 7021 49181 7055 49215
rect 7665 49181 7699 49215
rect 8217 49181 8251 49215
rect 4997 49113 5031 49147
rect 6469 49045 6503 49079
rect 7113 49045 7147 49079
rect 7481 49045 7515 49079
rect 8401 49045 8435 49079
rect 5089 48841 5123 48875
rect 5457 48841 5491 48875
rect 5825 48841 5859 48875
rect 7021 48773 7055 48807
rect 5273 48705 5307 48739
rect 5917 48637 5951 48671
rect 6009 48637 6043 48671
rect 6745 48637 6779 48671
rect 8493 48501 8527 48535
rect 7573 48297 7607 48331
rect 5457 48229 5491 48263
rect 6009 48161 6043 48195
rect 7021 48161 7055 48195
rect 5365 48093 5399 48127
rect 5825 48093 5859 48127
rect 7113 48093 7147 48127
rect 7205 48093 7239 48127
rect 5181 47957 5215 47991
rect 5917 47957 5951 47991
rect 6653 47753 6687 47787
rect 4721 47685 4755 47719
rect 7021 47685 7055 47719
rect 6469 47617 6503 47651
rect 4445 47549 4479 47583
rect 6745 47549 6779 47583
rect 6193 47413 6227 47447
rect 8493 47413 8527 47447
rect 6837 47209 6871 47243
rect 8401 47209 8435 47243
rect 6009 47073 6043 47107
rect 7297 47073 7331 47107
rect 7389 47073 7423 47107
rect 5825 47005 5859 47039
rect 6285 47005 6319 47039
rect 7205 47005 7239 47039
rect 8217 47005 8251 47039
rect 6653 46937 6687 46971
rect 5457 46869 5491 46903
rect 5917 46869 5951 46903
rect 7205 46529 7239 46563
rect 8217 46529 8251 46563
rect 4445 46461 4479 46495
rect 4721 46461 4755 46495
rect 6193 46461 6227 46495
rect 7297 46461 7331 46495
rect 7389 46461 7423 46495
rect 6837 46325 6871 46359
rect 8401 46325 8435 46359
rect 5181 46121 5215 46155
rect 8493 46121 8527 46155
rect 6101 45985 6135 46019
rect 5365 45917 5399 45951
rect 5917 45917 5951 45951
rect 6469 45917 6503 45951
rect 6745 45917 6779 45951
rect 7021 45849 7055 45883
rect 5549 45781 5583 45815
rect 6009 45781 6043 45815
rect 6653 45781 6687 45815
rect 6101 45577 6135 45611
rect 7297 45577 7331 45611
rect 7389 45509 7423 45543
rect 7757 45441 7791 45475
rect 4353 45373 4387 45407
rect 4629 45373 4663 45407
rect 7573 45373 7607 45407
rect 7941 45373 7975 45407
rect 6929 45237 6963 45271
rect 5273 45033 5307 45067
rect 8493 45033 8527 45067
rect 5457 44829 5491 44863
rect 6745 44829 6779 44863
rect 7021 44761 7055 44795
rect 7021 44489 7055 44523
rect 8401 44489 8435 44523
rect 5365 44353 5399 44387
rect 7205 44353 7239 44387
rect 8217 44353 8251 44387
rect 5181 44149 5215 44183
rect 6653 43945 6687 43979
rect 5181 43809 5215 43843
rect 4905 43741 4939 43775
rect 8493 43741 8527 43775
rect 8309 43605 8343 43639
rect 5365 43401 5399 43435
rect 5825 43401 5859 43435
rect 6745 43401 6779 43435
rect 5733 43265 5767 43299
rect 6929 43265 6963 43299
rect 7297 43265 7331 43299
rect 6009 43197 6043 43231
rect 6469 43197 6503 43231
rect 7113 43061 7147 43095
rect 6824 42857 6858 42891
rect 6561 42721 6595 42755
rect 4721 42653 4755 42687
rect 4997 42585 5031 42619
rect 6469 42517 6503 42551
rect 8309 42517 8343 42551
rect 5273 42313 5307 42347
rect 7297 42313 7331 42347
rect 7665 42313 7699 42347
rect 8033 42313 8067 42347
rect 5825 42245 5859 42279
rect 6009 42245 6043 42279
rect 6837 42245 6871 42279
rect 6929 42245 6963 42279
rect 8125 42245 8159 42279
rect 5457 42177 5491 42211
rect 5641 42177 5675 42211
rect 7481 42177 7515 42211
rect 6745 42109 6779 42143
rect 7849 42109 7883 42143
rect 8493 41973 8527 42007
rect 6561 41769 6595 41803
rect 5825 41565 5859 41599
rect 6469 41565 6503 41599
rect 7481 41565 7515 41599
rect 8217 41565 8251 41599
rect 6193 41497 6227 41531
rect 8033 41497 8067 41531
rect 7389 41429 7423 41463
rect 6193 41225 6227 41259
rect 4445 41089 4479 41123
rect 6469 41089 6503 41123
rect 8217 41089 8251 41123
rect 4721 41021 4755 41055
rect 6653 40885 6687 40919
rect 8401 40885 8435 40919
rect 4629 40681 4663 40715
rect 4813 40477 4847 40511
rect 6653 40477 6687 40511
rect 6745 40477 6779 40511
rect 7021 40409 7055 40443
rect 5365 40341 5399 40375
rect 8493 40341 8527 40375
rect 5273 40137 5307 40171
rect 5733 40137 5767 40171
rect 6745 40137 6779 40171
rect 7113 40137 7147 40171
rect 5641 40069 5675 40103
rect 6377 40001 6411 40035
rect 5917 39933 5951 39967
rect 7205 39933 7239 39967
rect 7389 39933 7423 39967
rect 6561 39797 6595 39831
rect 4721 39389 4755 39423
rect 6745 39389 6779 39423
rect 4997 39321 5031 39355
rect 7021 39321 7055 39355
rect 6469 39253 6503 39287
rect 8493 39253 8527 39287
rect 5181 39049 5215 39083
rect 5457 39049 5491 39083
rect 7481 39049 7515 39083
rect 7573 39049 7607 39083
rect 8401 39049 8435 39083
rect 5825 38981 5859 39015
rect 5365 38913 5399 38947
rect 5917 38913 5951 38947
rect 7021 38913 7055 38947
rect 7113 38913 7147 38947
rect 7757 38913 7791 38947
rect 8217 38913 8251 38947
rect 6101 38845 6135 38879
rect 6929 38845 6963 38879
rect 6745 38437 6779 38471
rect 4629 38301 4663 38335
rect 8217 38301 8251 38335
rect 4905 38233 4939 38267
rect 6561 38233 6595 38267
rect 6377 38165 6411 38199
rect 8401 38165 8435 38199
rect 5089 37961 5123 37995
rect 5457 37961 5491 37995
rect 5825 37961 5859 37995
rect 6653 37961 6687 37995
rect 7021 37893 7055 37927
rect 5273 37825 5307 37859
rect 6469 37825 6503 37859
rect 5917 37757 5951 37791
rect 6101 37757 6135 37791
rect 6745 37757 6779 37791
rect 8493 37621 8527 37655
rect 6745 37417 6779 37451
rect 6009 37281 6043 37315
rect 7297 37281 7331 37315
rect 5273 37213 5307 37247
rect 7113 37213 7147 37247
rect 5733 37145 5767 37179
rect 7205 37145 7239 37179
rect 5089 37077 5123 37111
rect 5365 37077 5399 37111
rect 5825 37077 5859 37111
rect 6193 36873 6227 36907
rect 6653 36873 6687 36907
rect 4721 36805 4755 36839
rect 7021 36805 7055 36839
rect 6469 36737 6503 36771
rect 4445 36669 4479 36703
rect 6745 36669 6779 36703
rect 8493 36533 8527 36567
rect 6653 36329 6687 36363
rect 8401 36329 8435 36363
rect 7113 36193 7147 36227
rect 7205 36193 7239 36227
rect 7021 36125 7055 36159
rect 8217 36125 8251 36159
rect 5825 35785 5859 35819
rect 5273 35649 5307 35683
rect 8217 35649 8251 35683
rect 5917 35581 5951 35615
rect 6101 35581 6135 35615
rect 5457 35513 5491 35547
rect 5089 35445 5123 35479
rect 8401 35445 8435 35479
rect 6377 35241 6411 35275
rect 4905 35105 4939 35139
rect 4629 35037 4663 35071
rect 6469 35037 6503 35071
rect 6745 35037 6779 35071
rect 7021 34969 7055 35003
rect 6653 34901 6687 34935
rect 8493 34901 8527 34935
rect 4629 34629 4663 34663
rect 5825 34561 5859 34595
rect 6837 34561 6871 34595
rect 5365 34493 5399 34527
rect 7573 34493 7607 34527
rect 5641 34357 5675 34391
rect 5076 34153 5110 34187
rect 6745 34017 6779 34051
rect 4813 33949 4847 33983
rect 7021 33881 7055 33915
rect 6561 33813 6595 33847
rect 8493 33813 8527 33847
rect 5457 33609 5491 33643
rect 5825 33609 5859 33643
rect 6745 33609 6779 33643
rect 7113 33609 7147 33643
rect 7941 33609 7975 33643
rect 5917 33541 5951 33575
rect 8033 33541 8067 33575
rect 7205 33473 7239 33507
rect 6101 33405 6135 33439
rect 7389 33405 7423 33439
rect 8125 33405 8159 33439
rect 7573 33269 7607 33303
rect 7021 33065 7055 33099
rect 7573 33065 7607 33099
rect 7205 32861 7239 32895
rect 7665 32861 7699 32895
rect 7941 32793 7975 32827
rect 8217 32725 8251 32759
rect 6653 32521 6687 32555
rect 7021 32453 7055 32487
rect 6469 32385 6503 32419
rect 4445 32317 4479 32351
rect 4721 32317 4755 32351
rect 6745 32317 6779 32351
rect 6193 32181 6227 32215
rect 8493 32181 8527 32215
rect 5089 31977 5123 32011
rect 6745 31977 6779 32011
rect 5549 31909 5583 31943
rect 6101 31841 6135 31875
rect 7205 31841 7239 31875
rect 7389 31841 7423 31875
rect 5273 31773 5307 31807
rect 7113 31773 7147 31807
rect 5457 31705 5491 31739
rect 5917 31705 5951 31739
rect 6009 31637 6043 31671
rect 6653 31433 6687 31467
rect 7021 31365 7055 31399
rect 6469 31297 6503 31331
rect 6745 31229 6779 31263
rect 8493 31093 8527 31127
rect 6745 30889 6779 30923
rect 7941 30889 7975 30923
rect 8401 30889 8435 30923
rect 4813 30753 4847 30787
rect 7205 30753 7239 30787
rect 7389 30753 7423 30787
rect 7113 30685 7147 30719
rect 8217 30685 8251 30719
rect 5089 30617 5123 30651
rect 7665 30617 7699 30651
rect 6561 30549 6595 30583
rect 5181 30345 5215 30379
rect 6745 30277 6779 30311
rect 5365 30209 5399 30243
rect 8217 30209 8251 30243
rect 6837 30141 6871 30175
rect 6929 30141 6963 30175
rect 6377 30073 6411 30107
rect 8401 30005 8435 30039
rect 6101 29665 6135 29699
rect 6009 29597 6043 29631
rect 6469 29597 6503 29631
rect 6745 29597 6779 29631
rect 7021 29529 7055 29563
rect 5549 29461 5583 29495
rect 5917 29461 5951 29495
rect 6653 29461 6687 29495
rect 8493 29461 8527 29495
rect 5457 29257 5491 29291
rect 6837 29257 6871 29291
rect 7205 29257 7239 29291
rect 5825 29189 5859 29223
rect 7297 29189 7331 29223
rect 5089 29121 5123 29155
rect 5365 29121 5399 29155
rect 5917 29121 5951 29155
rect 6101 29053 6135 29087
rect 7481 29053 7515 29087
rect 4905 28917 4939 28951
rect 5181 28917 5215 28951
rect 4813 28577 4847 28611
rect 5089 28577 5123 28611
rect 6745 28509 6779 28543
rect 7021 28441 7055 28475
rect 6561 28373 6595 28407
rect 8493 28373 8527 28407
rect 6193 28169 6227 28203
rect 7665 28169 7699 28203
rect 8401 28169 8435 28203
rect 7113 28101 7147 28135
rect 7205 28101 7239 28135
rect 4445 28033 4479 28067
rect 7849 28033 7883 28067
rect 8217 28033 8251 28067
rect 4721 27965 4755 27999
rect 7021 27965 7055 27999
rect 7573 27897 7607 27931
rect 8217 27421 8251 27455
rect 8493 27421 8527 27455
rect 8033 27285 8067 27319
rect 8309 27285 8343 27319
rect 7665 27013 7699 27047
rect 7757 26945 7791 26979
rect 8401 26945 8435 26979
rect 6929 26877 6963 26911
rect 7481 26877 7515 26911
rect 8125 26809 8159 26843
rect 6377 26741 6411 26775
rect 8217 26741 8251 26775
rect 4340 26537 4374 26571
rect 5825 26537 5859 26571
rect 7757 26537 7791 26571
rect 4077 26401 4111 26435
rect 5917 26401 5951 26435
rect 7665 26401 7699 26435
rect 8309 26401 8343 26435
rect 6193 26265 6227 26299
rect 6377 25993 6411 26027
rect 5733 25925 5767 25959
rect 8125 25925 8159 25959
rect 6561 25857 6595 25891
rect 6193 25789 6227 25823
rect 8401 25789 8435 25823
rect 6101 25721 6135 25755
rect 6653 25653 6687 25687
rect 7021 25313 7055 25347
rect 8217 25313 8251 25347
rect 8309 25313 8343 25347
rect 6929 25245 6963 25279
rect 7665 25177 7699 25211
rect 8125 25177 8159 25211
rect 6745 25109 6779 25143
rect 7757 25109 7791 25143
rect 6561 24769 6595 24803
rect 6837 24701 6871 24735
rect 8309 24565 8343 24599
rect 7389 24361 7423 24395
rect 8309 24225 8343 24259
rect 7297 24157 7331 24191
rect 8217 24089 8251 24123
rect 7757 24021 7791 24055
rect 8125 24021 8159 24055
rect 7849 23817 7883 23851
rect 6469 23681 6503 23715
rect 6837 23681 6871 23715
rect 8401 23681 8435 23715
rect 7205 23613 7239 23647
rect 7021 23545 7055 23579
rect 6653 23477 6687 23511
rect 7757 23477 7791 23511
rect 8309 23273 8343 23307
rect 6561 23069 6595 23103
rect 6837 23001 6871 23035
rect 7757 22729 7791 22763
rect 8125 22729 8159 22763
rect 8217 22661 8251 22695
rect 6929 22593 6963 22627
rect 7205 22593 7239 22627
rect 7481 22593 7515 22627
rect 8309 22525 8343 22559
rect 7665 22457 7699 22491
rect 7113 22389 7147 22423
rect 7389 22389 7423 22423
rect 8309 22049 8343 22083
rect 8033 21913 8067 21947
rect 6561 21845 6595 21879
rect 6929 21641 6963 21675
rect 8217 21641 8251 21675
rect 6745 21505 6779 21539
rect 7021 21505 7055 21539
rect 7665 21505 7699 21539
rect 8125 21505 8159 21539
rect 8309 21437 8343 21471
rect 7757 21301 7791 21335
rect 6561 20961 6595 20995
rect 6837 20825 6871 20859
rect 8309 20757 8343 20791
rect 7205 20553 7239 20587
rect 7389 20417 7423 20451
rect 7481 20417 7515 20451
rect 8125 20417 8159 20451
rect 8217 20349 8251 20383
rect 8309 20349 8343 20383
rect 7665 20281 7699 20315
rect 7757 20213 7791 20247
rect 7849 20009 7883 20043
rect 6837 19941 6871 19975
rect 8401 19873 8435 19907
rect 6561 19805 6595 19839
rect 7021 19805 7055 19839
rect 7205 19805 7239 19839
rect 6745 19669 6779 19703
rect 7757 19669 7791 19703
rect 8309 19465 8343 19499
rect 6837 19397 6871 19431
rect 6561 19329 6595 19363
rect 8217 18785 8251 18819
rect 8309 18785 8343 18819
rect 7389 18717 7423 18751
rect 8125 18717 8159 18751
rect 7205 18581 7239 18615
rect 7757 18581 7791 18615
rect 6837 18309 6871 18343
rect 6561 18241 6595 18275
rect 8309 18037 8343 18071
rect 7297 17765 7331 17799
rect 7665 17765 7699 17799
rect 8217 17697 8251 17731
rect 8309 17697 8343 17731
rect 7113 17629 7147 17663
rect 7481 17561 7515 17595
rect 7757 17493 7791 17527
rect 8125 17493 8159 17527
rect 7849 17289 7883 17323
rect 6561 17153 6595 17187
rect 7021 17153 7055 17187
rect 8401 17153 8435 17187
rect 7205 17085 7239 17119
rect 6837 17017 6871 17051
rect 6745 16949 6779 16983
rect 7757 16949 7791 16983
rect 8309 16745 8343 16779
rect 6561 16609 6595 16643
rect 6837 16609 6871 16643
rect 7757 16201 7791 16235
rect 8125 16201 8159 16235
rect 7205 16065 7239 16099
rect 8217 15997 8251 16031
rect 8309 15997 8343 16031
rect 7389 15861 7423 15895
rect 8033 15521 8067 15555
rect 8309 15453 8343 15487
rect 6561 15317 6595 15351
rect 7297 15045 7331 15079
rect 8033 15045 8067 15079
rect 6653 14977 6687 15011
rect 8493 14977 8527 15011
rect 7205 14773 7239 14807
rect 8309 14773 8343 14807
rect 7297 14501 7331 14535
rect 8217 14433 8251 14467
rect 8309 14433 8343 14467
rect 6837 14365 6871 14399
rect 7113 14365 7147 14399
rect 8125 14365 8159 14399
rect 6101 14297 6135 14331
rect 7573 14297 7607 14331
rect 6929 14229 6963 14263
rect 7757 14229 7791 14263
rect 6837 13957 6871 13991
rect 6561 13889 6595 13923
rect 8309 13821 8343 13855
rect 6653 13481 6687 13515
rect 7757 13413 7791 13447
rect 7113 13345 7147 13379
rect 8217 13345 8251 13379
rect 8401 13345 8435 13379
rect 6469 13277 6503 13311
rect 6929 13277 6963 13311
rect 7665 13209 7699 13243
rect 8125 13209 8159 13243
rect 6745 13141 6779 13175
rect 6837 12869 6871 12903
rect 6561 12801 6595 12835
rect 8309 12597 8343 12631
rect 8309 12257 8343 12291
rect 7481 12189 7515 12223
rect 8217 12121 8251 12155
rect 7665 12053 7699 12087
rect 7757 12053 7791 12087
rect 8125 12053 8159 12087
rect 6745 11849 6779 11883
rect 7849 11849 7883 11883
rect 6561 11713 6595 11747
rect 7021 11713 7055 11747
rect 8401 11713 8435 11747
rect 7205 11645 7239 11679
rect 6837 11509 6871 11543
rect 7757 11509 7791 11543
rect 8309 11305 8343 11339
rect 6561 11169 6595 11203
rect 6837 11169 6871 11203
rect 7757 10761 7791 10795
rect 8125 10761 8159 10795
rect 7389 10625 7423 10659
rect 8217 10557 8251 10591
rect 8401 10557 8435 10591
rect 7205 10421 7239 10455
rect 6561 10081 6595 10115
rect 6837 10081 6871 10115
rect 8309 9877 8343 9911
rect 7481 9537 7515 9571
rect 8125 9537 8159 9571
rect 8217 9469 8251 9503
rect 8401 9469 8435 9503
rect 7665 9401 7699 9435
rect 7757 9333 7791 9367
rect 6745 9129 6779 9163
rect 7849 9129 7883 9163
rect 8401 8993 8435 9027
rect 6561 8925 6595 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 6837 8789 6871 8823
rect 7757 8789 7791 8823
rect 8309 8585 8343 8619
rect 6561 8449 6595 8483
rect 6009 8381 6043 8415
rect 6837 8381 6871 8415
rect 5457 8245 5491 8279
rect 5181 7905 5215 7939
rect 6929 7905 6963 7939
rect 7573 7905 7607 7939
rect 8217 7905 8251 7939
rect 8309 7905 8343 7939
rect 4629 7837 4663 7871
rect 5089 7837 5123 7871
rect 8125 7837 8159 7871
rect 4721 7769 4755 7803
rect 4905 7769 4939 7803
rect 5457 7769 5491 7803
rect 4445 7701 4479 7735
rect 7021 7701 7055 7735
rect 7757 7701 7791 7735
rect 5917 7497 5951 7531
rect 4261 7429 4295 7463
rect 3709 7361 3743 7395
rect 6101 7361 6135 7395
rect 6377 7361 6411 7395
rect 6653 7361 6687 7395
rect 3985 7293 4019 7327
rect 5733 7293 5767 7327
rect 6929 7293 6963 7327
rect 6561 7225 6595 7259
rect 3893 7157 3927 7191
rect 8401 7157 8435 7191
rect 4058 6953 4092 6987
rect 6009 6953 6043 6987
rect 7757 6953 7791 6987
rect 6193 6885 6227 6919
rect 7573 6817 7607 6851
rect 8309 6817 8343 6851
rect 3801 6749 3835 6783
rect 7297 6749 7331 6783
rect 6469 6681 6503 6715
rect 5549 6613 5583 6647
rect 8125 6613 8159 6647
rect 8217 6613 8251 6647
rect 7389 6409 7423 6443
rect 7849 6409 7883 6443
rect 7665 6341 7699 6375
rect 8401 6273 8435 6307
rect 8309 5865 8343 5899
rect 8493 5661 8527 5695
rect 1869 3009 1903 3043
rect 2329 3009 2363 3043
rect 2421 3009 2455 3043
rect 1685 2805 1719 2839
rect 2145 2805 2179 2839
rect 7573 2601 7607 2635
rect 7941 2601 7975 2635
rect 1869 2465 1903 2499
rect 6653 2465 6687 2499
rect 4445 2397 4479 2431
rect 6377 2397 6411 2431
rect 8125 2397 8159 2431
rect 7665 2329 7699 2363
rect 8493 2329 8527 2363
rect 4169 2261 4203 2295
<< metal1 >>
rect 1104 77818 8832 77840
rect 1104 77766 2350 77818
rect 2402 77766 2414 77818
rect 2466 77766 2478 77818
rect 2530 77766 2542 77818
rect 2594 77766 2606 77818
rect 2658 77766 7350 77818
rect 7402 77766 7414 77818
rect 7466 77766 7478 77818
rect 7530 77766 7542 77818
rect 7594 77766 7606 77818
rect 7658 77766 8832 77818
rect 1104 77744 8832 77766
rect 2682 77460 2688 77512
rect 2740 77460 2746 77512
rect 2869 77435 2927 77441
rect 2869 77401 2881 77435
rect 2915 77432 2927 77435
rect 5534 77432 5540 77444
rect 2915 77404 5540 77432
rect 2915 77401 2927 77404
rect 2869 77395 2927 77401
rect 5534 77392 5540 77404
rect 5592 77392 5598 77444
rect 1104 77274 8832 77296
rect 1104 77222 3010 77274
rect 3062 77222 3074 77274
rect 3126 77222 3138 77274
rect 3190 77222 3202 77274
rect 3254 77222 3266 77274
rect 3318 77222 8010 77274
rect 8062 77222 8074 77274
rect 8126 77222 8138 77274
rect 8190 77222 8202 77274
rect 8254 77222 8266 77274
rect 8318 77222 8832 77274
rect 1104 77200 8832 77222
rect 1104 76730 8832 76752
rect 1104 76678 2350 76730
rect 2402 76678 2414 76730
rect 2466 76678 2478 76730
rect 2530 76678 2542 76730
rect 2594 76678 2606 76730
rect 2658 76678 7350 76730
rect 7402 76678 7414 76730
rect 7466 76678 7478 76730
rect 7530 76678 7542 76730
rect 7594 76678 7606 76730
rect 7658 76678 8832 76730
rect 1104 76656 8832 76678
rect 1104 76186 8832 76208
rect 1104 76134 3010 76186
rect 3062 76134 3074 76186
rect 3126 76134 3138 76186
rect 3190 76134 3202 76186
rect 3254 76134 3266 76186
rect 3318 76134 8010 76186
rect 8062 76134 8074 76186
rect 8126 76134 8138 76186
rect 8190 76134 8202 76186
rect 8254 76134 8266 76186
rect 8318 76134 8832 76186
rect 1104 76112 8832 76134
rect 1104 75642 8832 75664
rect 1104 75590 2350 75642
rect 2402 75590 2414 75642
rect 2466 75590 2478 75642
rect 2530 75590 2542 75642
rect 2594 75590 2606 75642
rect 2658 75590 7350 75642
rect 7402 75590 7414 75642
rect 7466 75590 7478 75642
rect 7530 75590 7542 75642
rect 7594 75590 7606 75642
rect 7658 75590 8832 75642
rect 1104 75568 8832 75590
rect 1104 75098 8832 75120
rect 1104 75046 3010 75098
rect 3062 75046 3074 75098
rect 3126 75046 3138 75098
rect 3190 75046 3202 75098
rect 3254 75046 3266 75098
rect 3318 75046 8010 75098
rect 8062 75046 8074 75098
rect 8126 75046 8138 75098
rect 8190 75046 8202 75098
rect 8254 75046 8266 75098
rect 8318 75046 8832 75098
rect 1104 75024 8832 75046
rect 1104 74554 8832 74576
rect 1104 74502 2350 74554
rect 2402 74502 2414 74554
rect 2466 74502 2478 74554
rect 2530 74502 2542 74554
rect 2594 74502 2606 74554
rect 2658 74502 7350 74554
rect 7402 74502 7414 74554
rect 7466 74502 7478 74554
rect 7530 74502 7542 74554
rect 7594 74502 7606 74554
rect 7658 74502 8832 74554
rect 1104 74480 8832 74502
rect 7926 74196 7932 74248
rect 7984 74236 7990 74248
rect 8205 74239 8263 74245
rect 8205 74236 8217 74239
rect 7984 74208 8217 74236
rect 7984 74196 7990 74208
rect 8205 74205 8217 74208
rect 8251 74205 8263 74239
rect 8205 74199 8263 74205
rect 8386 74060 8392 74112
rect 8444 74060 8450 74112
rect 1104 74010 8832 74032
rect 1104 73958 3010 74010
rect 3062 73958 3074 74010
rect 3126 73958 3138 74010
rect 3190 73958 3202 74010
rect 3254 73958 3266 74010
rect 3318 73958 8010 74010
rect 8062 73958 8074 74010
rect 8126 73958 8138 74010
rect 8190 73958 8202 74010
rect 8254 73958 8266 74010
rect 8318 73958 8832 74010
rect 1104 73936 8832 73958
rect 7742 73788 7748 73840
rect 7800 73788 7806 73840
rect 5534 73720 5540 73772
rect 5592 73760 5598 73772
rect 6362 73760 6368 73772
rect 5592 73732 6368 73760
rect 5592 73720 5598 73732
rect 6362 73720 6368 73732
rect 6420 73720 6426 73772
rect 6730 73652 6736 73704
rect 6788 73652 6794 73704
rect 7006 73652 7012 73704
rect 7064 73652 7070 73704
rect 6549 73559 6607 73565
rect 6549 73525 6561 73559
rect 6595 73556 6607 73559
rect 6638 73556 6644 73568
rect 6595 73528 6644 73556
rect 6595 73525 6607 73528
rect 6549 73519 6607 73525
rect 6638 73516 6644 73528
rect 6696 73516 6702 73568
rect 8018 73516 8024 73568
rect 8076 73556 8082 73568
rect 8481 73559 8539 73565
rect 8481 73556 8493 73559
rect 8076 73528 8493 73556
rect 8076 73516 8082 73528
rect 8481 73525 8493 73528
rect 8527 73525 8539 73559
rect 8481 73519 8539 73525
rect 1104 73466 8832 73488
rect 1104 73414 2350 73466
rect 2402 73414 2414 73466
rect 2466 73414 2478 73466
rect 2530 73414 2542 73466
rect 2594 73414 2606 73466
rect 2658 73414 7350 73466
rect 7402 73414 7414 73466
rect 7466 73414 7478 73466
rect 7530 73414 7542 73466
rect 7594 73414 7606 73466
rect 7658 73414 8832 73466
rect 1104 73392 8832 73414
rect 7006 73312 7012 73364
rect 7064 73352 7070 73364
rect 7745 73355 7803 73361
rect 7745 73352 7757 73355
rect 7064 73324 7757 73352
rect 7064 73312 7070 73324
rect 7745 73321 7757 73324
rect 7791 73321 7803 73355
rect 7745 73315 7803 73321
rect 7834 73284 7840 73296
rect 7116 73256 7840 73284
rect 7116 73225 7144 73256
rect 7834 73244 7840 73256
rect 7892 73244 7898 73296
rect 7101 73219 7159 73225
rect 7101 73185 7113 73219
rect 7147 73185 7159 73219
rect 8018 73216 8024 73228
rect 7101 73179 7159 73185
rect 7300 73188 8024 73216
rect 5074 73108 5080 73160
rect 5132 73108 5138 73160
rect 7300 73157 7328 73188
rect 8018 73176 8024 73188
rect 8076 73176 8082 73228
rect 7285 73151 7343 73157
rect 7285 73117 7297 73151
rect 7331 73117 7343 73151
rect 7929 73151 7987 73157
rect 7929 73148 7941 73151
rect 7285 73111 7343 73117
rect 7484 73120 7941 73148
rect 5350 73040 5356 73092
rect 5408 73040 5414 73092
rect 6638 73080 6644 73092
rect 6578 73052 6644 73080
rect 6638 73040 6644 73052
rect 6696 73040 6702 73092
rect 6822 72972 6828 73024
rect 6880 73012 6886 73024
rect 7193 73015 7251 73021
rect 7193 73012 7205 73015
rect 6880 72984 7205 73012
rect 6880 72972 6886 72984
rect 7193 72981 7205 72984
rect 7239 72981 7251 73015
rect 7484 73012 7512 73120
rect 7929 73117 7941 73120
rect 7975 73117 7987 73151
rect 7929 73111 7987 73117
rect 8018 73040 8024 73092
rect 8076 73080 8082 73092
rect 8113 73083 8171 73089
rect 8113 73080 8125 73083
rect 8076 73052 8125 73080
rect 8076 73040 8082 73052
rect 8113 73049 8125 73052
rect 8159 73049 8171 73083
rect 8113 73043 8171 73049
rect 7653 73015 7711 73021
rect 7653 73012 7665 73015
rect 7484 72984 7665 73012
rect 7193 72975 7251 72981
rect 7653 72981 7665 72984
rect 7699 72981 7711 73015
rect 7653 72975 7711 72981
rect 7742 72972 7748 73024
rect 7800 73012 7806 73024
rect 8205 73015 8263 73021
rect 8205 73012 8217 73015
rect 7800 72984 8217 73012
rect 7800 72972 7806 72984
rect 8205 72981 8217 72984
rect 8251 72981 8263 73015
rect 8205 72975 8263 72981
rect 1104 72922 8832 72944
rect 1104 72870 3010 72922
rect 3062 72870 3074 72922
rect 3126 72870 3138 72922
rect 3190 72870 3202 72922
rect 3254 72870 3266 72922
rect 3318 72870 8010 72922
rect 8062 72870 8074 72922
rect 8126 72870 8138 72922
rect 8190 72870 8202 72922
rect 8254 72870 8266 72922
rect 8318 72870 8832 72922
rect 1104 72848 8832 72870
rect 5350 72768 5356 72820
rect 5408 72808 5414 72820
rect 5445 72811 5503 72817
rect 5445 72808 5457 72811
rect 5408 72780 5457 72808
rect 5408 72768 5414 72780
rect 5445 72777 5457 72780
rect 5491 72777 5503 72811
rect 5445 72771 5503 72777
rect 6365 72811 6423 72817
rect 6365 72777 6377 72811
rect 6411 72777 6423 72811
rect 6365 72771 6423 72777
rect 5629 72675 5687 72681
rect 5629 72641 5641 72675
rect 5675 72672 5687 72675
rect 6380 72672 6408 72771
rect 6638 72768 6644 72820
rect 6696 72808 6702 72820
rect 7926 72808 7932 72820
rect 6696 72780 7932 72808
rect 6696 72768 6702 72780
rect 7926 72768 7932 72780
rect 7984 72768 7990 72820
rect 5675 72644 6408 72672
rect 5675 72641 5687 72644
rect 5629 72635 5687 72641
rect 6638 72632 6644 72684
rect 6696 72672 6702 72684
rect 6733 72675 6791 72681
rect 6733 72672 6745 72675
rect 6696 72644 6745 72672
rect 6696 72632 6702 72644
rect 6733 72641 6745 72644
rect 6779 72641 6791 72675
rect 6733 72635 6791 72641
rect 7006 72632 7012 72684
rect 7064 72672 7070 72684
rect 7377 72675 7435 72681
rect 7377 72672 7389 72675
rect 7064 72644 7389 72672
rect 7064 72632 7070 72644
rect 7377 72641 7389 72644
rect 7423 72641 7435 72675
rect 7377 72635 7435 72641
rect 6822 72564 6828 72616
rect 6880 72564 6886 72616
rect 6917 72607 6975 72613
rect 6917 72573 6929 72607
rect 6963 72573 6975 72607
rect 6917 72567 6975 72573
rect 6454 72428 6460 72480
rect 6512 72468 6518 72480
rect 6932 72468 6960 72567
rect 6512 72440 6960 72468
rect 6512 72428 6518 72440
rect 7098 72428 7104 72480
rect 7156 72468 7162 72480
rect 7193 72471 7251 72477
rect 7193 72468 7205 72471
rect 7156 72440 7205 72468
rect 7156 72428 7162 72440
rect 7193 72437 7205 72440
rect 7239 72437 7251 72471
rect 7193 72431 7251 72437
rect 1104 72378 8832 72400
rect 1104 72326 2350 72378
rect 2402 72326 2414 72378
rect 2466 72326 2478 72378
rect 2530 72326 2542 72378
rect 2594 72326 2606 72378
rect 2658 72326 7350 72378
rect 7402 72326 7414 72378
rect 7466 72326 7478 72378
rect 7530 72326 7542 72378
rect 7594 72326 7606 72378
rect 7658 72326 8832 72378
rect 1104 72304 8832 72326
rect 4430 72088 4436 72140
rect 4488 72128 4494 72140
rect 4801 72131 4859 72137
rect 4801 72128 4813 72131
rect 4488 72100 4813 72128
rect 4488 72088 4494 72100
rect 4801 72097 4813 72100
rect 4847 72128 4859 72131
rect 5074 72128 5080 72140
rect 4847 72100 5080 72128
rect 4847 72097 4859 72100
rect 4801 72091 4859 72097
rect 5074 72088 5080 72100
rect 5132 72088 5138 72140
rect 6730 72088 6736 72140
rect 6788 72088 6794 72140
rect 7009 72131 7067 72137
rect 7009 72097 7021 72131
rect 7055 72128 7067 72131
rect 7098 72128 7104 72140
rect 7055 72100 7104 72128
rect 7055 72097 7067 72100
rect 7009 72091 7067 72097
rect 7098 72088 7104 72100
rect 7156 72088 7162 72140
rect 6546 72060 6552 72072
rect 6210 72046 6552 72060
rect 6196 72032 6552 72046
rect 5074 71952 5080 72004
rect 5132 71952 5138 72004
rect 5810 71884 5816 71936
rect 5868 71924 5874 71936
rect 6196 71924 6224 72032
rect 6546 72020 6552 72032
rect 6604 72020 6610 72072
rect 7098 71952 7104 72004
rect 7156 71992 7162 72004
rect 7156 71964 7498 71992
rect 7156 71952 7162 71964
rect 5868 71896 6224 71924
rect 5868 71884 5874 71896
rect 6546 71884 6552 71936
rect 6604 71884 6610 71936
rect 7392 71924 7420 71964
rect 7742 71924 7748 71936
rect 7392 71896 7748 71924
rect 7742 71884 7748 71896
rect 7800 71884 7806 71936
rect 7926 71884 7932 71936
rect 7984 71924 7990 71936
rect 8481 71927 8539 71933
rect 8481 71924 8493 71927
rect 7984 71896 8493 71924
rect 7984 71884 7990 71896
rect 8481 71893 8493 71896
rect 8527 71893 8539 71927
rect 8481 71887 8539 71893
rect 1104 71834 8832 71856
rect 1104 71782 3010 71834
rect 3062 71782 3074 71834
rect 3126 71782 3138 71834
rect 3190 71782 3202 71834
rect 3254 71782 3266 71834
rect 3318 71782 8010 71834
rect 8062 71782 8074 71834
rect 8126 71782 8138 71834
rect 8190 71782 8202 71834
rect 8254 71782 8266 71834
rect 8318 71782 8832 71834
rect 1104 71760 8832 71782
rect 5074 71680 5080 71732
rect 5132 71720 5138 71732
rect 5261 71723 5319 71729
rect 5261 71720 5273 71723
rect 5132 71692 5273 71720
rect 5132 71680 5138 71692
rect 5261 71689 5273 71692
rect 5307 71689 5319 71723
rect 5261 71683 5319 71689
rect 6365 71723 6423 71729
rect 6365 71689 6377 71723
rect 6411 71689 6423 71723
rect 6365 71683 6423 71689
rect 6733 71723 6791 71729
rect 6733 71689 6745 71723
rect 6779 71720 6791 71723
rect 6822 71720 6828 71732
rect 6779 71692 6828 71720
rect 6779 71689 6791 71692
rect 6733 71683 6791 71689
rect 5445 71587 5503 71593
rect 5445 71553 5457 71587
rect 5491 71584 5503 71587
rect 6380 71584 6408 71683
rect 6822 71680 6828 71692
rect 6880 71680 6886 71732
rect 7006 71680 7012 71732
rect 7064 71720 7070 71732
rect 7193 71723 7251 71729
rect 7193 71720 7205 71723
rect 7064 71692 7205 71720
rect 7064 71680 7070 71692
rect 7193 71689 7205 71692
rect 7239 71689 7251 71723
rect 7193 71683 7251 71689
rect 8389 71723 8447 71729
rect 8389 71689 8401 71723
rect 8435 71720 8447 71723
rect 8478 71720 8484 71732
rect 8435 71692 8484 71720
rect 8435 71689 8447 71692
rect 8389 71683 8447 71689
rect 8478 71680 8484 71692
rect 8536 71680 8542 71732
rect 7561 71655 7619 71661
rect 7561 71621 7573 71655
rect 7607 71652 7619 71655
rect 7926 71652 7932 71664
rect 7607 71624 7932 71652
rect 7607 71621 7619 71624
rect 7561 71615 7619 71621
rect 7926 71612 7932 71624
rect 7984 71652 7990 71664
rect 8113 71655 8171 71661
rect 8113 71652 8125 71655
rect 7984 71624 8125 71652
rect 7984 71612 7990 71624
rect 8113 71621 8125 71624
rect 8159 71621 8171 71655
rect 8113 71615 8171 71621
rect 7653 71587 7711 71593
rect 7653 71584 7665 71587
rect 5491 71556 6408 71584
rect 6840 71556 7665 71584
rect 5491 71553 5503 71556
rect 5445 71547 5503 71553
rect 5902 71476 5908 71528
rect 5960 71516 5966 71528
rect 6546 71516 6552 71528
rect 5960 71488 6552 71516
rect 5960 71476 5966 71488
rect 6546 71476 6552 71488
rect 6604 71516 6610 71528
rect 6840 71525 6868 71556
rect 7653 71553 7665 71556
rect 7699 71553 7711 71587
rect 7653 71547 7711 71553
rect 6825 71519 6883 71525
rect 6825 71516 6837 71519
rect 6604 71488 6837 71516
rect 6604 71476 6610 71488
rect 6825 71485 6837 71488
rect 6871 71485 6883 71519
rect 6825 71479 6883 71485
rect 6917 71519 6975 71525
rect 6917 71485 6929 71519
rect 6963 71485 6975 71519
rect 6917 71479 6975 71485
rect 6454 71448 6460 71460
rect 6104 71420 6460 71448
rect 6104 71392 6132 71420
rect 6454 71408 6460 71420
rect 6512 71448 6518 71460
rect 6932 71448 6960 71479
rect 7834 71476 7840 71528
rect 7892 71476 7898 71528
rect 6512 71420 6960 71448
rect 6512 71408 6518 71420
rect 6086 71340 6092 71392
rect 6144 71340 6150 71392
rect 1104 71290 8832 71312
rect 1104 71238 2350 71290
rect 2402 71238 2414 71290
rect 2466 71238 2478 71290
rect 2530 71238 2542 71290
rect 2594 71238 2606 71290
rect 2658 71238 7350 71290
rect 7402 71238 7414 71290
rect 7466 71238 7478 71290
rect 7530 71238 7542 71290
rect 7594 71238 7606 71290
rect 7658 71238 8832 71290
rect 1104 71216 8832 71238
rect 6086 71000 6092 71052
rect 6144 71000 6150 71052
rect 5353 70975 5411 70981
rect 5353 70941 5365 70975
rect 5399 70972 5411 70975
rect 5399 70944 5580 70972
rect 5399 70941 5411 70944
rect 5353 70935 5411 70941
rect 4982 70796 4988 70848
rect 5040 70836 5046 70848
rect 5552 70845 5580 70944
rect 5902 70932 5908 70984
rect 5960 70932 5966 70984
rect 6914 70932 6920 70984
rect 6972 70972 6978 70984
rect 7193 70975 7251 70981
rect 7193 70972 7205 70975
rect 6972 70944 7205 70972
rect 6972 70932 6978 70944
rect 7193 70941 7205 70944
rect 7239 70941 7251 70975
rect 7193 70935 7251 70941
rect 7926 70932 7932 70984
rect 7984 70972 7990 70984
rect 8205 70975 8263 70981
rect 8205 70972 8217 70975
rect 7984 70944 8217 70972
rect 7984 70932 7990 70944
rect 8205 70941 8217 70944
rect 8251 70941 8263 70975
rect 8205 70935 8263 70941
rect 5169 70839 5227 70845
rect 5169 70836 5181 70839
rect 5040 70808 5181 70836
rect 5040 70796 5046 70808
rect 5169 70805 5181 70808
rect 5215 70805 5227 70839
rect 5169 70799 5227 70805
rect 5537 70839 5595 70845
rect 5537 70805 5549 70839
rect 5583 70805 5595 70839
rect 5537 70799 5595 70805
rect 5997 70839 6055 70845
rect 5997 70805 6009 70839
rect 6043 70836 6055 70839
rect 6178 70836 6184 70848
rect 6043 70808 6184 70836
rect 6043 70805 6055 70808
rect 5997 70799 6055 70805
rect 6178 70796 6184 70808
rect 6236 70796 6242 70848
rect 7006 70796 7012 70848
rect 7064 70796 7070 70848
rect 8386 70796 8392 70848
rect 8444 70796 8450 70848
rect 1104 70746 8832 70768
rect 1104 70694 3010 70746
rect 3062 70694 3074 70746
rect 3126 70694 3138 70746
rect 3190 70694 3202 70746
rect 3254 70694 3266 70746
rect 3318 70694 8010 70746
rect 8062 70694 8074 70746
rect 8126 70694 8138 70746
rect 8190 70694 8202 70746
rect 8254 70694 8266 70746
rect 8318 70694 8832 70746
rect 1104 70672 8832 70694
rect 4709 70567 4767 70573
rect 4709 70533 4721 70567
rect 4755 70564 4767 70567
rect 4982 70564 4988 70576
rect 4755 70536 4988 70564
rect 4755 70533 4767 70536
rect 4709 70527 4767 70533
rect 4982 70524 4988 70536
rect 5040 70524 5046 70576
rect 7006 70524 7012 70576
rect 7064 70524 7070 70576
rect 7098 70524 7104 70576
rect 7156 70564 7162 70576
rect 7156 70536 7498 70564
rect 7156 70524 7162 70536
rect 4430 70456 4436 70508
rect 4488 70456 4494 70508
rect 5810 70456 5816 70508
rect 5868 70496 5874 70508
rect 5868 70468 6684 70496
rect 5868 70456 5874 70468
rect 6178 70388 6184 70440
rect 6236 70388 6242 70440
rect 6656 70428 6684 70468
rect 6730 70456 6736 70508
rect 6788 70456 6794 70508
rect 7006 70428 7012 70440
rect 6656 70400 7012 70428
rect 7006 70388 7012 70400
rect 7064 70388 7070 70440
rect 8481 70431 8539 70437
rect 8481 70428 8493 70431
rect 8036 70400 8493 70428
rect 8036 70372 8064 70400
rect 8481 70397 8493 70400
rect 8527 70397 8539 70431
rect 8481 70391 8539 70397
rect 8018 70320 8024 70372
rect 8076 70320 8082 70372
rect 1104 70202 8832 70224
rect 1104 70150 2350 70202
rect 2402 70150 2414 70202
rect 2466 70150 2478 70202
rect 2530 70150 2542 70202
rect 2594 70150 2606 70202
rect 2658 70150 7350 70202
rect 7402 70150 7414 70202
rect 7466 70150 7478 70202
rect 7530 70150 7542 70202
rect 7594 70150 7606 70202
rect 7658 70150 8832 70202
rect 1104 70128 8832 70150
rect 6914 70048 6920 70100
rect 6972 70048 6978 70100
rect 7561 69955 7619 69961
rect 7561 69921 7573 69955
rect 7607 69952 7619 69955
rect 7834 69952 7840 69964
rect 7607 69924 7840 69952
rect 7607 69921 7619 69924
rect 7561 69915 7619 69921
rect 7834 69912 7840 69924
rect 7892 69912 7898 69964
rect 7285 69887 7343 69893
rect 7285 69853 7297 69887
rect 7331 69884 7343 69887
rect 7926 69884 7932 69896
rect 7331 69856 7932 69884
rect 7331 69853 7343 69856
rect 7285 69847 7343 69853
rect 7926 69844 7932 69856
rect 7984 69844 7990 69896
rect 5902 69708 5908 69760
rect 5960 69748 5966 69760
rect 6178 69748 6184 69760
rect 5960 69720 6184 69748
rect 5960 69708 5966 69720
rect 6178 69708 6184 69720
rect 6236 69748 6242 69760
rect 7377 69751 7435 69757
rect 7377 69748 7389 69751
rect 6236 69720 7389 69748
rect 6236 69708 6242 69720
rect 7377 69717 7389 69720
rect 7423 69717 7435 69751
rect 7377 69711 7435 69717
rect 1104 69658 8832 69680
rect 1104 69606 3010 69658
rect 3062 69606 3074 69658
rect 3126 69606 3138 69658
rect 3190 69606 3202 69658
rect 3254 69606 3266 69658
rect 3318 69606 8010 69658
rect 8062 69606 8074 69658
rect 8126 69606 8138 69658
rect 8190 69606 8202 69658
rect 8254 69606 8266 69658
rect 8318 69606 8832 69658
rect 1104 69584 8832 69606
rect 4430 69368 4436 69420
rect 4488 69368 4494 69420
rect 7098 69408 7104 69420
rect 5842 69380 7104 69408
rect 7098 69368 7104 69380
rect 7156 69368 7162 69420
rect 7193 69411 7251 69417
rect 7193 69377 7205 69411
rect 7239 69408 7251 69411
rect 8205 69411 8263 69417
rect 8205 69408 8217 69411
rect 7239 69380 8217 69408
rect 7239 69377 7251 69380
rect 7193 69371 7251 69377
rect 8205 69377 8217 69380
rect 8251 69408 8263 69411
rect 8478 69408 8484 69420
rect 8251 69380 8484 69408
rect 8251 69377 8263 69380
rect 8205 69371 8263 69377
rect 8478 69368 8484 69380
rect 8536 69368 8542 69420
rect 4706 69300 4712 69352
rect 4764 69300 4770 69352
rect 5994 69300 6000 69352
rect 6052 69340 6058 69352
rect 6181 69343 6239 69349
rect 6181 69340 6193 69343
rect 6052 69312 6193 69340
rect 6052 69300 6058 69312
rect 6181 69309 6193 69312
rect 6227 69340 6239 69343
rect 7285 69343 7343 69349
rect 7285 69340 7297 69343
rect 6227 69312 7297 69340
rect 6227 69309 6239 69312
rect 6181 69303 6239 69309
rect 7285 69309 7297 69312
rect 7331 69309 7343 69343
rect 7285 69303 7343 69309
rect 7469 69343 7527 69349
rect 7469 69309 7481 69343
rect 7515 69340 7527 69343
rect 7834 69340 7840 69352
rect 7515 69312 7840 69340
rect 7515 69309 7527 69312
rect 7469 69303 7527 69309
rect 7834 69300 7840 69312
rect 7892 69300 7898 69352
rect 6638 69164 6644 69216
rect 6696 69204 6702 69216
rect 6825 69207 6883 69213
rect 6825 69204 6837 69207
rect 6696 69176 6837 69204
rect 6696 69164 6702 69176
rect 6825 69173 6837 69176
rect 6871 69173 6883 69207
rect 6825 69167 6883 69173
rect 8386 69164 8392 69216
rect 8444 69164 8450 69216
rect 1104 69114 8832 69136
rect 1104 69062 2350 69114
rect 2402 69062 2414 69114
rect 2466 69062 2478 69114
rect 2530 69062 2542 69114
rect 2594 69062 2606 69114
rect 2658 69062 7350 69114
rect 7402 69062 7414 69114
rect 7466 69062 7478 69114
rect 7530 69062 7542 69114
rect 7594 69062 7606 69114
rect 7658 69062 8832 69114
rect 1104 69040 8832 69062
rect 4706 68960 4712 69012
rect 4764 69000 4770 69012
rect 5169 69003 5227 69009
rect 5169 69000 5181 69003
rect 4764 68972 5181 69000
rect 4764 68960 4770 68972
rect 5169 68969 5181 68972
rect 5215 68969 5227 69003
rect 5169 68963 5227 68969
rect 8478 68960 8484 69012
rect 8536 68960 8542 69012
rect 5994 68824 6000 68876
rect 6052 68824 6058 68876
rect 6181 68867 6239 68873
rect 6181 68833 6193 68867
rect 6227 68864 6239 68867
rect 6270 68864 6276 68876
rect 6227 68836 6276 68864
rect 6227 68833 6239 68836
rect 6181 68827 6239 68833
rect 6270 68824 6276 68836
rect 6328 68824 6334 68876
rect 5353 68799 5411 68805
rect 5353 68765 5365 68799
rect 5399 68796 5411 68799
rect 5399 68768 5580 68796
rect 5399 68765 5411 68768
rect 5353 68759 5411 68765
rect 5552 68669 5580 68768
rect 5902 68756 5908 68808
rect 5960 68756 5966 68808
rect 6457 68799 6515 68805
rect 6457 68765 6469 68799
rect 6503 68796 6515 68799
rect 6638 68796 6644 68808
rect 6503 68768 6644 68796
rect 6503 68765 6515 68768
rect 6457 68759 6515 68765
rect 6638 68756 6644 68768
rect 6696 68756 6702 68808
rect 6730 68756 6736 68808
rect 6788 68756 6794 68808
rect 7009 68731 7067 68737
rect 7009 68728 7021 68731
rect 6656 68700 7021 68728
rect 6656 68669 6684 68700
rect 7009 68697 7021 68700
rect 7055 68697 7067 68731
rect 7009 68691 7067 68697
rect 7098 68688 7104 68740
rect 7156 68728 7162 68740
rect 7156 68700 7498 68728
rect 7156 68688 7162 68700
rect 5537 68663 5595 68669
rect 5537 68629 5549 68663
rect 5583 68629 5595 68663
rect 5537 68623 5595 68629
rect 6641 68663 6699 68669
rect 6641 68629 6653 68663
rect 6687 68629 6699 68663
rect 6641 68623 6699 68629
rect 1104 68570 8832 68592
rect 1104 68518 3010 68570
rect 3062 68518 3074 68570
rect 3126 68518 3138 68570
rect 3190 68518 3202 68570
rect 3254 68518 3266 68570
rect 3318 68518 8010 68570
rect 8062 68518 8074 68570
rect 8126 68518 8138 68570
rect 8190 68518 8202 68570
rect 8254 68518 8266 68570
rect 8318 68518 8832 68570
rect 1104 68496 8832 68518
rect 5445 68459 5503 68465
rect 5445 68425 5457 68459
rect 5491 68425 5503 68459
rect 5445 68419 5503 68425
rect 5813 68459 5871 68465
rect 5813 68425 5825 68459
rect 5859 68456 5871 68459
rect 5994 68456 6000 68468
rect 5859 68428 6000 68456
rect 5859 68425 5871 68428
rect 5813 68419 5871 68425
rect 5353 68323 5411 68329
rect 5353 68289 5365 68323
rect 5399 68320 5411 68323
rect 5460 68320 5488 68419
rect 5994 68416 6000 68428
rect 6052 68416 6058 68468
rect 5399 68292 5488 68320
rect 5905 68323 5963 68329
rect 5399 68289 5411 68292
rect 5353 68283 5411 68289
rect 5905 68289 5917 68323
rect 5951 68320 5963 68323
rect 6546 68320 6552 68332
rect 5951 68292 6552 68320
rect 5951 68289 5963 68292
rect 5905 68283 5963 68289
rect 6546 68280 6552 68292
rect 6604 68320 6610 68332
rect 7101 68323 7159 68329
rect 7101 68320 7113 68323
rect 6604 68292 7113 68320
rect 6604 68280 6610 68292
rect 7101 68289 7113 68292
rect 7147 68289 7159 68323
rect 7101 68283 7159 68289
rect 7193 68323 7251 68329
rect 7193 68289 7205 68323
rect 7239 68320 7251 68323
rect 8205 68323 8263 68329
rect 8205 68320 8217 68323
rect 7239 68292 8217 68320
rect 7239 68289 7251 68292
rect 7193 68283 7251 68289
rect 8205 68289 8217 68292
rect 8251 68320 8263 68323
rect 8251 68292 8800 68320
rect 8251 68289 8263 68292
rect 8205 68283 8263 68289
rect 6089 68255 6147 68261
rect 6089 68221 6101 68255
rect 6135 68252 6147 68255
rect 6822 68252 6828 68264
rect 6135 68224 6828 68252
rect 6135 68221 6147 68224
rect 6089 68215 6147 68221
rect 6822 68212 6828 68224
rect 6880 68212 6886 68264
rect 7009 68255 7067 68261
rect 7009 68221 7021 68255
rect 7055 68252 7067 68255
rect 7834 68252 7840 68264
rect 7055 68224 7840 68252
rect 7055 68221 7067 68224
rect 7009 68215 7067 68221
rect 7834 68212 7840 68224
rect 7892 68212 7898 68264
rect 5166 68076 5172 68128
rect 5224 68076 5230 68128
rect 7561 68119 7619 68125
rect 7561 68085 7573 68119
rect 7607 68116 7619 68119
rect 7742 68116 7748 68128
rect 7607 68088 7748 68116
rect 7607 68085 7619 68088
rect 7561 68079 7619 68085
rect 7742 68076 7748 68088
rect 7800 68076 7806 68128
rect 8386 68076 8392 68128
rect 8444 68076 8450 68128
rect 8772 68116 8800 68292
rect 8772 68088 8892 68116
rect 1104 68026 8832 68048
rect 1104 67974 2350 68026
rect 2402 67974 2414 68026
rect 2466 67974 2478 68026
rect 2530 67974 2542 68026
rect 2594 67974 2606 68026
rect 2658 67974 7350 68026
rect 7402 67974 7414 68026
rect 7466 67974 7478 68026
rect 7530 67974 7542 68026
rect 7594 67974 7606 68026
rect 7658 67974 8832 68026
rect 1104 67952 8832 67974
rect 6546 67872 6552 67924
rect 6604 67872 6610 67924
rect 8481 67915 8539 67921
rect 8481 67881 8493 67915
rect 8527 67912 8539 67915
rect 8864 67912 8892 68088
rect 8527 67884 8892 67912
rect 8527 67881 8539 67884
rect 8481 67875 8539 67881
rect 4430 67736 4436 67788
rect 4488 67776 4494 67788
rect 4801 67779 4859 67785
rect 4801 67776 4813 67779
rect 4488 67748 4813 67776
rect 4488 67736 4494 67748
rect 4801 67745 4813 67748
rect 4847 67745 4859 67779
rect 4801 67739 4859 67745
rect 5077 67779 5135 67785
rect 5077 67745 5089 67779
rect 5123 67776 5135 67779
rect 5166 67776 5172 67788
rect 5123 67748 5172 67776
rect 5123 67745 5135 67748
rect 5077 67739 5135 67745
rect 5166 67736 5172 67748
rect 5224 67736 5230 67788
rect 7006 67736 7012 67788
rect 7064 67776 7070 67788
rect 7650 67776 7656 67788
rect 7064 67748 7656 67776
rect 7064 67736 7070 67748
rect 7650 67736 7656 67748
rect 7708 67736 7714 67788
rect 6730 67668 6736 67720
rect 6788 67668 6794 67720
rect 6302 67612 6592 67640
rect 6086 67532 6092 67584
rect 6144 67572 6150 67584
rect 6564 67572 6592 67612
rect 7006 67600 7012 67652
rect 7064 67600 7070 67652
rect 7098 67600 7104 67652
rect 7156 67640 7162 67652
rect 7156 67612 7498 67640
rect 7156 67600 7162 67612
rect 7116 67572 7144 67600
rect 6144 67544 7144 67572
rect 6144 67532 6150 67544
rect 1104 67482 8832 67504
rect 1104 67430 3010 67482
rect 3062 67430 3074 67482
rect 3126 67430 3138 67482
rect 3190 67430 3202 67482
rect 3254 67430 3266 67482
rect 3318 67430 8010 67482
rect 8062 67430 8074 67482
rect 8126 67430 8138 67482
rect 8190 67430 8202 67482
rect 8254 67430 8266 67482
rect 8318 67430 8832 67482
rect 1104 67408 8832 67430
rect 6546 67328 6552 67380
rect 6604 67368 6610 67380
rect 6733 67371 6791 67377
rect 6733 67368 6745 67371
rect 6604 67340 6745 67368
rect 6604 67328 6610 67340
rect 6733 67337 6745 67340
rect 6779 67337 6791 67371
rect 6733 67331 6791 67337
rect 7006 67328 7012 67380
rect 7064 67368 7070 67380
rect 7193 67371 7251 67377
rect 7193 67368 7205 67371
rect 7064 67340 7205 67368
rect 7064 67328 7070 67340
rect 7193 67337 7205 67340
rect 7239 67337 7251 67371
rect 7193 67331 7251 67337
rect 7742 67328 7748 67380
rect 7800 67328 7806 67380
rect 6825 67303 6883 67309
rect 6825 67269 6837 67303
rect 6871 67300 6883 67303
rect 6914 67300 6920 67312
rect 6871 67272 6920 67300
rect 6871 67269 6883 67272
rect 6825 67263 6883 67269
rect 6914 67260 6920 67272
rect 6972 67260 6978 67312
rect 7377 67235 7435 67241
rect 7377 67201 7389 67235
rect 7423 67232 7435 67235
rect 7760 67232 7788 67328
rect 7423 67204 7788 67232
rect 8205 67235 8263 67241
rect 7423 67201 7435 67204
rect 7377 67195 7435 67201
rect 8205 67201 8217 67235
rect 8251 67232 8263 67235
rect 8478 67232 8484 67244
rect 8251 67204 8484 67232
rect 8251 67201 8263 67204
rect 8205 67195 8263 67201
rect 8478 67192 8484 67204
rect 8536 67192 8542 67244
rect 6822 67124 6828 67176
rect 6880 67164 6886 67176
rect 6917 67167 6975 67173
rect 6917 67164 6929 67167
rect 6880 67136 6929 67164
rect 6880 67124 6886 67136
rect 6917 67133 6929 67136
rect 6963 67133 6975 67167
rect 6917 67127 6975 67133
rect 6362 66988 6368 67040
rect 6420 66988 6426 67040
rect 8386 66988 8392 67040
rect 8444 66988 8450 67040
rect 1104 66938 8832 66960
rect 1104 66886 2350 66938
rect 2402 66886 2414 66938
rect 2466 66886 2478 66938
rect 2530 66886 2542 66938
rect 2594 66886 2606 66938
rect 2658 66886 7350 66938
rect 7402 66886 7414 66938
rect 7466 66886 7478 66938
rect 7530 66886 7542 66938
rect 7594 66886 7606 66938
rect 7658 66886 8832 66938
rect 1104 66864 8832 66886
rect 6549 66827 6607 66833
rect 6549 66793 6561 66827
rect 6595 66824 6607 66827
rect 6914 66824 6920 66836
rect 6595 66796 6920 66824
rect 6595 66793 6607 66796
rect 6549 66787 6607 66793
rect 6914 66784 6920 66796
rect 6972 66784 6978 66836
rect 4430 66648 4436 66700
rect 4488 66688 4494 66700
rect 4801 66691 4859 66697
rect 4801 66688 4813 66691
rect 4488 66660 4813 66688
rect 4488 66648 4494 66660
rect 4801 66657 4813 66660
rect 4847 66657 4859 66691
rect 6932 66688 6960 66784
rect 8113 66691 8171 66697
rect 8113 66688 8125 66691
rect 6932 66660 8125 66688
rect 4801 66651 4859 66657
rect 8113 66657 8125 66660
rect 8159 66657 8171 66691
rect 8113 66651 8171 66657
rect 8205 66691 8263 66697
rect 8205 66657 8217 66691
rect 8251 66657 8263 66691
rect 8205 66651 8263 66657
rect 6086 66580 6092 66632
rect 6144 66620 6150 66632
rect 7006 66620 7012 66632
rect 6144 66592 7012 66620
rect 6144 66580 6150 66592
rect 7006 66580 7012 66592
rect 7064 66580 7070 66632
rect 7098 66580 7104 66632
rect 7156 66620 7162 66632
rect 7834 66620 7840 66632
rect 7156 66592 7840 66620
rect 7156 66580 7162 66592
rect 7834 66580 7840 66592
rect 7892 66620 7898 66632
rect 8220 66620 8248 66651
rect 7892 66592 8248 66620
rect 7892 66580 7898 66592
rect 5074 66512 5080 66564
rect 5132 66512 5138 66564
rect 6641 66555 6699 66561
rect 6641 66552 6653 66555
rect 6380 66524 6653 66552
rect 5718 66444 5724 66496
rect 5776 66484 5782 66496
rect 6380 66484 6408 66524
rect 6641 66521 6653 66524
rect 6687 66521 6699 66555
rect 6641 66515 6699 66521
rect 6730 66512 6736 66564
rect 6788 66552 6794 66564
rect 7377 66555 7435 66561
rect 7377 66552 7389 66555
rect 6788 66524 7389 66552
rect 6788 66512 6794 66524
rect 7377 66521 7389 66524
rect 7423 66521 7435 66555
rect 7377 66515 7435 66521
rect 8021 66555 8079 66561
rect 8021 66521 8033 66555
rect 8067 66552 8079 66555
rect 8067 66524 8524 66552
rect 8067 66521 8079 66524
rect 8021 66515 8079 66521
rect 8496 66496 8524 66524
rect 5776 66456 6408 66484
rect 5776 66444 5782 66456
rect 7650 66444 7656 66496
rect 7708 66444 7714 66496
rect 8478 66444 8484 66496
rect 8536 66444 8542 66496
rect 1104 66394 8832 66416
rect 1104 66342 3010 66394
rect 3062 66342 3074 66394
rect 3126 66342 3138 66394
rect 3190 66342 3202 66394
rect 3254 66342 3266 66394
rect 3318 66342 8010 66394
rect 8062 66342 8074 66394
rect 8126 66342 8138 66394
rect 8190 66342 8202 66394
rect 8254 66342 8266 66394
rect 8318 66342 8832 66394
rect 1104 66320 8832 66342
rect 5074 66240 5080 66292
rect 5132 66280 5138 66292
rect 5261 66283 5319 66289
rect 5261 66280 5273 66283
rect 5132 66252 5273 66280
rect 5132 66240 5138 66252
rect 5261 66249 5273 66252
rect 5307 66249 5319 66283
rect 5261 66243 5319 66249
rect 6362 66240 6368 66292
rect 6420 66240 6426 66292
rect 7650 66280 7656 66292
rect 6932 66252 7656 66280
rect 5445 66147 5503 66153
rect 5445 66113 5457 66147
rect 5491 66144 5503 66147
rect 6380 66144 6408 66240
rect 6932 66212 6960 66252
rect 7650 66240 7656 66252
rect 7708 66240 7714 66292
rect 8478 66240 8484 66292
rect 8536 66240 8542 66292
rect 6472 66184 6960 66212
rect 6472 66153 6500 66184
rect 7006 66172 7012 66224
rect 7064 66212 7070 66224
rect 7064 66184 7498 66212
rect 7064 66172 7070 66184
rect 5491 66116 6408 66144
rect 6457 66147 6515 66153
rect 5491 66113 5503 66116
rect 5445 66107 5503 66113
rect 6457 66113 6469 66147
rect 6503 66113 6515 66147
rect 6457 66107 6515 66113
rect 6730 66036 6736 66088
rect 6788 66036 6794 66088
rect 7009 66079 7067 66085
rect 7009 66076 7021 66079
rect 6840 66048 7021 66076
rect 6641 66011 6699 66017
rect 6641 65977 6653 66011
rect 6687 66008 6699 66011
rect 6840 66008 6868 66048
rect 7009 66045 7021 66048
rect 7055 66045 7067 66079
rect 7009 66039 7067 66045
rect 6687 65980 6868 66008
rect 6687 65977 6699 65980
rect 6641 65971 6699 65977
rect 1104 65850 8832 65872
rect 1104 65798 2350 65850
rect 2402 65798 2414 65850
rect 2466 65798 2478 65850
rect 2530 65798 2542 65850
rect 2594 65798 2606 65850
rect 2658 65798 7350 65850
rect 7402 65798 7414 65850
rect 7466 65798 7478 65850
rect 7530 65798 7542 65850
rect 7594 65798 7606 65850
rect 7658 65798 8832 65850
rect 1104 65776 8832 65798
rect 4430 65560 4436 65612
rect 4488 65600 4494 65612
rect 4801 65603 4859 65609
rect 4801 65600 4813 65603
rect 4488 65572 4813 65600
rect 4488 65560 4494 65572
rect 4801 65569 4813 65572
rect 4847 65569 4859 65603
rect 4801 65563 4859 65569
rect 5810 65560 5816 65612
rect 5868 65600 5874 65612
rect 6822 65600 6828 65612
rect 5868 65572 6828 65600
rect 5868 65560 5874 65572
rect 6822 65560 6828 65572
rect 6880 65600 6886 65612
rect 7469 65603 7527 65609
rect 7469 65600 7481 65603
rect 6880 65572 7481 65600
rect 6880 65560 6886 65572
rect 7469 65569 7481 65572
rect 7515 65569 7527 65603
rect 7469 65563 7527 65569
rect 6086 65492 6092 65544
rect 6144 65532 6150 65544
rect 6144 65504 6210 65532
rect 6144 65492 6150 65504
rect 6914 65492 6920 65544
rect 6972 65532 6978 65544
rect 7285 65535 7343 65541
rect 7285 65532 7297 65535
rect 6972 65504 7297 65532
rect 6972 65492 6978 65504
rect 7285 65501 7297 65504
rect 7331 65501 7343 65535
rect 7285 65495 7343 65501
rect 7926 65492 7932 65544
rect 7984 65532 7990 65544
rect 8205 65535 8263 65541
rect 8205 65532 8217 65535
rect 7984 65504 8217 65532
rect 7984 65492 7990 65504
rect 8205 65501 8217 65504
rect 8251 65501 8263 65535
rect 8205 65495 8263 65501
rect 5074 65424 5080 65476
rect 5132 65424 5138 65476
rect 6825 65467 6883 65473
rect 6825 65433 6837 65467
rect 6871 65464 6883 65467
rect 6871 65436 7420 65464
rect 6871 65433 6883 65436
rect 6825 65427 6883 65433
rect 6914 65356 6920 65408
rect 6972 65356 6978 65408
rect 7392 65405 7420 65436
rect 7377 65399 7435 65405
rect 7377 65365 7389 65399
rect 7423 65396 7435 65399
rect 7742 65396 7748 65408
rect 7423 65368 7748 65396
rect 7423 65365 7435 65368
rect 7377 65359 7435 65365
rect 7742 65356 7748 65368
rect 7800 65356 7806 65408
rect 8386 65356 8392 65408
rect 8444 65356 8450 65408
rect 1104 65306 8832 65328
rect 1104 65254 3010 65306
rect 3062 65254 3074 65306
rect 3126 65254 3138 65306
rect 3190 65254 3202 65306
rect 3254 65254 3266 65306
rect 3318 65254 8010 65306
rect 8062 65254 8074 65306
rect 8126 65254 8138 65306
rect 8190 65254 8202 65306
rect 8254 65254 8266 65306
rect 8318 65254 8832 65306
rect 1104 65232 8832 65254
rect 5074 65152 5080 65204
rect 5132 65192 5138 65204
rect 5629 65195 5687 65201
rect 5629 65192 5641 65195
rect 5132 65164 5641 65192
rect 5132 65152 5138 65164
rect 5629 65161 5641 65164
rect 5675 65161 5687 65195
rect 5629 65155 5687 65161
rect 6914 65152 6920 65204
rect 6972 65152 6978 65204
rect 4430 65084 4436 65136
rect 4488 65124 4494 65136
rect 4709 65127 4767 65133
rect 4709 65124 4721 65127
rect 4488 65096 4721 65124
rect 4488 65084 4494 65096
rect 4709 65093 4721 65096
rect 4755 65093 4767 65127
rect 6932 65124 6960 65152
rect 4709 65087 4767 65093
rect 5828 65096 6960 65124
rect 5534 65016 5540 65068
rect 5592 65016 5598 65068
rect 5828 65065 5856 65096
rect 7834 65084 7840 65136
rect 7892 65124 7898 65136
rect 8113 65127 8171 65133
rect 8113 65124 8125 65127
rect 7892 65096 8125 65124
rect 7892 65084 7898 65096
rect 8113 65093 8125 65096
rect 8159 65093 8171 65127
rect 8113 65087 8171 65093
rect 5813 65059 5871 65065
rect 5813 65025 5825 65059
rect 5859 65025 5871 65059
rect 5813 65019 5871 65025
rect 6825 65059 6883 65065
rect 6825 65025 6837 65059
rect 6871 65056 6883 65059
rect 7098 65056 7104 65068
rect 6871 65028 7104 65056
rect 6871 65025 6883 65028
rect 6825 65019 6883 65025
rect 7098 65016 7104 65028
rect 7156 65016 7162 65068
rect 7006 64812 7012 64864
rect 7064 64812 7070 64864
rect 8202 64812 8208 64864
rect 8260 64812 8266 64864
rect 1104 64762 8832 64784
rect 1104 64710 2350 64762
rect 2402 64710 2414 64762
rect 2466 64710 2478 64762
rect 2530 64710 2542 64762
rect 2594 64710 2606 64762
rect 2658 64710 7350 64762
rect 7402 64710 7414 64762
rect 7466 64710 7478 64762
rect 7530 64710 7542 64762
rect 7594 64710 7606 64762
rect 7658 64710 8832 64762
rect 1104 64688 8832 64710
rect 7006 64472 7012 64524
rect 7064 64472 7070 64524
rect 7650 64472 7656 64524
rect 7708 64512 7714 64524
rect 8202 64512 8208 64524
rect 7708 64484 8208 64512
rect 7708 64472 7714 64484
rect 8202 64472 8208 64484
rect 8260 64472 8266 64524
rect 6454 64404 6460 64456
rect 6512 64404 6518 64456
rect 6730 64404 6736 64456
rect 6788 64404 6794 64456
rect 8220 64444 8248 64472
rect 8142 64416 8248 64444
rect 6638 64268 6644 64320
rect 6696 64268 6702 64320
rect 7926 64268 7932 64320
rect 7984 64308 7990 64320
rect 8481 64311 8539 64317
rect 8481 64308 8493 64311
rect 7984 64280 8493 64308
rect 7984 64268 7990 64280
rect 8481 64277 8493 64280
rect 8527 64277 8539 64311
rect 8481 64271 8539 64277
rect 1104 64218 8832 64240
rect 1104 64166 3010 64218
rect 3062 64166 3074 64218
rect 3126 64166 3138 64218
rect 3190 64166 3202 64218
rect 3254 64166 3266 64218
rect 3318 64166 8010 64218
rect 8062 64166 8074 64218
rect 8126 64166 8138 64218
rect 8190 64166 8202 64218
rect 8254 64166 8266 64218
rect 8318 64166 8832 64218
rect 1104 64144 8832 64166
rect 5261 64107 5319 64113
rect 5261 64073 5273 64107
rect 5307 64073 5319 64107
rect 5261 64067 5319 64073
rect 4985 63971 5043 63977
rect 4985 63937 4997 63971
rect 5031 63968 5043 63971
rect 5276 63968 5304 64067
rect 6638 64064 6644 64116
rect 6696 64064 6702 64116
rect 7006 64064 7012 64116
rect 7064 64104 7070 64116
rect 7650 64104 7656 64116
rect 7064 64076 7656 64104
rect 7064 64064 7070 64076
rect 7650 64064 7656 64076
rect 7708 64104 7714 64116
rect 7708 64076 7880 64104
rect 7708 64064 7714 64076
rect 6656 64036 6684 64064
rect 6733 64039 6791 64045
rect 6733 64036 6745 64039
rect 6656 64008 6745 64036
rect 6733 64005 6745 64008
rect 6779 64005 6791 64039
rect 6733 63999 6791 64005
rect 5031 63940 5304 63968
rect 5629 63971 5687 63977
rect 5031 63937 5043 63940
rect 4985 63931 5043 63937
rect 5629 63937 5641 63971
rect 5675 63968 5687 63971
rect 5902 63968 5908 63980
rect 5675 63940 5908 63968
rect 5675 63937 5687 63940
rect 5629 63931 5687 63937
rect 5902 63928 5908 63940
rect 5960 63928 5966 63980
rect 7852 63954 7880 64076
rect 5718 63860 5724 63912
rect 5776 63860 5782 63912
rect 5810 63860 5816 63912
rect 5868 63860 5874 63912
rect 6457 63903 6515 63909
rect 6457 63869 6469 63903
rect 6503 63869 6515 63903
rect 6457 63863 6515 63869
rect 4798 63724 4804 63776
rect 4856 63724 4862 63776
rect 6472 63764 6500 63863
rect 6730 63764 6736 63776
rect 6472 63736 6736 63764
rect 6730 63724 6736 63736
rect 6788 63724 6794 63776
rect 8202 63724 8208 63776
rect 8260 63724 8266 63776
rect 1104 63674 8832 63696
rect 1104 63622 2350 63674
rect 2402 63622 2414 63674
rect 2466 63622 2478 63674
rect 2530 63622 2542 63674
rect 2594 63622 2606 63674
rect 2658 63622 7350 63674
rect 7402 63622 7414 63674
rect 7466 63622 7478 63674
rect 7530 63622 7542 63674
rect 7594 63622 7606 63674
rect 7658 63622 8832 63674
rect 1104 63600 8832 63622
rect 4604 63563 4662 63569
rect 4604 63529 4616 63563
rect 4650 63560 4662 63563
rect 4798 63560 4804 63572
rect 4650 63532 4804 63560
rect 4650 63529 4662 63532
rect 4604 63523 4662 63529
rect 4798 63520 4804 63532
rect 4856 63520 4862 63572
rect 5718 63520 5724 63572
rect 5776 63560 5782 63572
rect 6089 63563 6147 63569
rect 6089 63560 6101 63563
rect 5776 63532 6101 63560
rect 5776 63520 5782 63532
rect 6089 63529 6101 63532
rect 6135 63529 6147 63563
rect 6089 63523 6147 63529
rect 6365 63563 6423 63569
rect 6365 63529 6377 63563
rect 6411 63560 6423 63563
rect 6454 63560 6460 63572
rect 6411 63532 6460 63560
rect 6411 63529 6423 63532
rect 6365 63523 6423 63529
rect 4338 63384 4344 63436
rect 4396 63384 4402 63436
rect 6104 63424 6132 63523
rect 6454 63520 6460 63532
rect 6512 63520 6518 63572
rect 7834 63520 7840 63572
rect 7892 63520 7898 63572
rect 8478 63560 8484 63572
rect 8404 63532 8484 63560
rect 7098 63452 7104 63504
rect 7156 63492 7162 63504
rect 7193 63495 7251 63501
rect 7193 63492 7205 63495
rect 7156 63464 7205 63492
rect 7156 63452 7162 63464
rect 7193 63461 7205 63464
rect 7239 63461 7251 63495
rect 7193 63455 7251 63461
rect 7282 63452 7288 63504
rect 7340 63492 7346 63504
rect 7852 63492 7880 63520
rect 8404 63501 8432 63532
rect 8478 63520 8484 63532
rect 8536 63520 8542 63572
rect 7340 63464 7880 63492
rect 8389 63495 8447 63501
rect 7340 63452 7346 63464
rect 8389 63461 8401 63495
rect 8435 63461 8447 63495
rect 8389 63455 8447 63461
rect 6825 63427 6883 63433
rect 6825 63424 6837 63427
rect 6104 63396 6837 63424
rect 6825 63393 6837 63396
rect 6871 63393 6883 63427
rect 6825 63387 6883 63393
rect 7009 63427 7067 63433
rect 7009 63393 7021 63427
rect 7055 63424 7067 63427
rect 7834 63424 7840 63436
rect 7055 63396 7840 63424
rect 7055 63393 7067 63396
rect 7009 63387 7067 63393
rect 7834 63384 7840 63396
rect 7892 63384 7898 63436
rect 6733 63359 6791 63365
rect 5750 63328 6316 63356
rect 5902 63248 5908 63300
rect 5960 63248 5966 63300
rect 6288 63288 6316 63328
rect 6733 63325 6745 63359
rect 6779 63356 6791 63359
rect 8113 63359 8171 63365
rect 8113 63356 8125 63359
rect 6779 63328 8125 63356
rect 6779 63325 6791 63328
rect 6733 63319 6791 63325
rect 8113 63325 8125 63328
rect 8159 63356 8171 63359
rect 8202 63356 8208 63368
rect 8159 63328 8208 63356
rect 8159 63325 8171 63328
rect 8113 63319 8171 63325
rect 8202 63316 8208 63328
rect 8260 63316 8266 63368
rect 7098 63288 7104 63300
rect 6288 63260 7104 63288
rect 7098 63248 7104 63260
rect 7156 63288 7162 63300
rect 7282 63288 7288 63300
rect 7156 63260 7288 63288
rect 7156 63248 7162 63260
rect 7282 63248 7288 63260
rect 7340 63248 7346 63300
rect 7561 63291 7619 63297
rect 7561 63257 7573 63291
rect 7607 63288 7619 63291
rect 7926 63288 7932 63300
rect 7607 63260 7932 63288
rect 7607 63257 7619 63260
rect 7561 63251 7619 63257
rect 7926 63248 7932 63260
rect 7984 63248 7990 63300
rect 5920 63220 5948 63248
rect 6638 63220 6644 63232
rect 5920 63192 6644 63220
rect 6638 63180 6644 63192
rect 6696 63220 6702 63232
rect 7653 63223 7711 63229
rect 7653 63220 7665 63223
rect 6696 63192 7665 63220
rect 6696 63180 6702 63192
rect 7653 63189 7665 63192
rect 7699 63189 7711 63223
rect 7653 63183 7711 63189
rect 1104 63130 8832 63152
rect 1104 63078 3010 63130
rect 3062 63078 3074 63130
rect 3126 63078 3138 63130
rect 3190 63078 3202 63130
rect 3254 63078 3266 63130
rect 3318 63078 8010 63130
rect 8062 63078 8074 63130
rect 8126 63078 8138 63130
rect 8190 63078 8202 63130
rect 8254 63078 8266 63130
rect 8318 63078 8832 63130
rect 1104 63056 8832 63078
rect 5537 63019 5595 63025
rect 5537 62985 5549 63019
rect 5583 63016 5595 63019
rect 5718 63016 5724 63028
rect 5583 62988 5724 63016
rect 5583 62985 5595 62988
rect 5537 62979 5595 62985
rect 5718 62976 5724 62988
rect 5776 62976 5782 63028
rect 4985 62883 5043 62889
rect 4985 62849 4997 62883
rect 5031 62880 5043 62883
rect 5629 62883 5687 62889
rect 5031 62852 5212 62880
rect 5031 62849 5043 62852
rect 4985 62843 5043 62849
rect 5184 62753 5212 62852
rect 5629 62849 5641 62883
rect 5675 62880 5687 62883
rect 5675 62852 6132 62880
rect 5675 62849 5687 62852
rect 5629 62843 5687 62849
rect 6104 62824 6132 62852
rect 8018 62840 8024 62892
rect 8076 62880 8082 62892
rect 8205 62883 8263 62889
rect 8205 62880 8217 62883
rect 8076 62852 8217 62880
rect 8076 62840 8082 62852
rect 8205 62849 8217 62852
rect 8251 62849 8263 62883
rect 8205 62843 8263 62849
rect 5813 62815 5871 62821
rect 5813 62781 5825 62815
rect 5859 62812 5871 62815
rect 5902 62812 5908 62824
rect 5859 62784 5908 62812
rect 5859 62781 5871 62784
rect 5813 62775 5871 62781
rect 5902 62772 5908 62784
rect 5960 62772 5966 62824
rect 6086 62772 6092 62824
rect 6144 62772 6150 62824
rect 5169 62747 5227 62753
rect 5169 62713 5181 62747
rect 5215 62713 5227 62747
rect 5169 62707 5227 62713
rect 4706 62636 4712 62688
rect 4764 62676 4770 62688
rect 4801 62679 4859 62685
rect 4801 62676 4813 62679
rect 4764 62648 4813 62676
rect 4764 62636 4770 62648
rect 4801 62645 4813 62648
rect 4847 62645 4859 62679
rect 4801 62639 4859 62645
rect 8386 62636 8392 62688
rect 8444 62636 8450 62688
rect 1104 62586 8832 62608
rect 1104 62534 2350 62586
rect 2402 62534 2414 62586
rect 2466 62534 2478 62586
rect 2530 62534 2542 62586
rect 2594 62534 2606 62586
rect 2658 62534 7350 62586
rect 7402 62534 7414 62586
rect 7466 62534 7478 62586
rect 7530 62534 7542 62586
rect 7594 62534 7606 62586
rect 7658 62534 8832 62586
rect 1104 62512 8832 62534
rect 7098 62472 7104 62484
rect 5736 62444 7104 62472
rect 4338 62296 4344 62348
rect 4396 62296 4402 62348
rect 4617 62339 4675 62345
rect 4617 62305 4629 62339
rect 4663 62336 4675 62339
rect 4706 62336 4712 62348
rect 4663 62308 4712 62336
rect 4663 62305 4675 62308
rect 4617 62299 4675 62305
rect 4706 62296 4712 62308
rect 4764 62296 4770 62348
rect 5736 62254 5764 62444
rect 7098 62432 7104 62444
rect 7156 62432 7162 62484
rect 7006 62296 7012 62348
rect 7064 62336 7070 62348
rect 7064 62308 8156 62336
rect 7064 62296 7070 62308
rect 6454 62228 6460 62280
rect 6512 62228 6518 62280
rect 6730 62228 6736 62280
rect 6788 62228 6794 62280
rect 8128 62254 8156 62308
rect 7009 62203 7067 62209
rect 7009 62169 7021 62203
rect 7055 62169 7067 62203
rect 7009 62163 7067 62169
rect 6086 62092 6092 62144
rect 6144 62092 6150 62144
rect 6641 62135 6699 62141
rect 6641 62101 6653 62135
rect 6687 62132 6699 62135
rect 7024 62132 7052 62163
rect 6687 62104 7052 62132
rect 6687 62101 6699 62104
rect 6641 62095 6699 62101
rect 7098 62092 7104 62144
rect 7156 62132 7162 62144
rect 8018 62132 8024 62144
rect 7156 62104 8024 62132
rect 7156 62092 7162 62104
rect 8018 62092 8024 62104
rect 8076 62132 8082 62144
rect 8481 62135 8539 62141
rect 8481 62132 8493 62135
rect 8076 62104 8493 62132
rect 8076 62092 8082 62104
rect 8481 62101 8493 62104
rect 8527 62101 8539 62135
rect 8481 62095 8539 62101
rect 1104 62042 8832 62064
rect 1104 61990 3010 62042
rect 3062 61990 3074 62042
rect 3126 61990 3138 62042
rect 3190 61990 3202 62042
rect 3254 61990 3266 62042
rect 3318 61990 8010 62042
rect 8062 61990 8074 62042
rect 8126 61990 8138 62042
rect 8190 61990 8202 62042
rect 8254 61990 8266 62042
rect 8318 61990 8832 62042
rect 1104 61968 8832 61990
rect 6454 61888 6460 61940
rect 6512 61928 6518 61940
rect 6733 61931 6791 61937
rect 6733 61928 6745 61931
rect 6512 61900 6745 61928
rect 6512 61888 6518 61900
rect 6733 61897 6745 61900
rect 6779 61897 6791 61931
rect 6733 61891 6791 61897
rect 7098 61888 7104 61940
rect 7156 61888 7162 61940
rect 6086 61820 6092 61872
rect 6144 61860 6150 61872
rect 7193 61863 7251 61869
rect 7193 61860 7205 61863
rect 6144 61832 7205 61860
rect 6144 61820 6150 61832
rect 7193 61829 7205 61832
rect 7239 61829 7251 61863
rect 7193 61823 7251 61829
rect 7377 61727 7435 61733
rect 7377 61693 7389 61727
rect 7423 61693 7435 61727
rect 7377 61687 7435 61693
rect 7098 61548 7104 61600
rect 7156 61588 7162 61600
rect 7392 61588 7420 61687
rect 7156 61560 7420 61588
rect 7156 61548 7162 61560
rect 1104 61498 8832 61520
rect 1104 61446 2350 61498
rect 2402 61446 2414 61498
rect 2466 61446 2478 61498
rect 2530 61446 2542 61498
rect 2594 61446 2606 61498
rect 2658 61446 7350 61498
rect 7402 61446 7414 61498
rect 7466 61446 7478 61498
rect 7530 61446 7542 61498
rect 7594 61446 7606 61498
rect 7658 61446 8832 61498
rect 1104 61424 8832 61446
rect 4338 61208 4344 61260
rect 4396 61248 4402 61260
rect 4433 61251 4491 61257
rect 4433 61248 4445 61251
rect 4396 61220 4445 61248
rect 4396 61208 4402 61220
rect 4433 61217 4445 61220
rect 4479 61217 4491 61251
rect 4433 61211 4491 61217
rect 6822 61140 6828 61192
rect 6880 61140 6886 61192
rect 7742 61140 7748 61192
rect 7800 61180 7806 61192
rect 8205 61183 8263 61189
rect 8205 61180 8217 61183
rect 7800 61152 8217 61180
rect 7800 61140 7806 61152
rect 8205 61149 8217 61152
rect 8251 61149 8263 61183
rect 8205 61143 8263 61149
rect 4706 61072 4712 61124
rect 4764 61072 4770 61124
rect 6914 61112 6920 61124
rect 5934 61084 6920 61112
rect 6914 61072 6920 61084
rect 6972 61072 6978 61124
rect 7469 61115 7527 61121
rect 7469 61081 7481 61115
rect 7515 61112 7527 61115
rect 7926 61112 7932 61124
rect 7515 61084 7932 61112
rect 7515 61081 7527 61084
rect 7469 61075 7527 61081
rect 7926 61072 7932 61084
rect 7984 61072 7990 61124
rect 5718 61004 5724 61056
rect 5776 61044 5782 61056
rect 6181 61047 6239 61053
rect 6181 61044 6193 61047
rect 5776 61016 6193 61044
rect 5776 61004 5782 61016
rect 6181 61013 6193 61016
rect 6227 61013 6239 61047
rect 6181 61007 6239 61013
rect 7006 61004 7012 61056
rect 7064 61004 7070 61056
rect 7098 61004 7104 61056
rect 7156 61044 7162 61056
rect 7374 61044 7380 61056
rect 7156 61016 7380 61044
rect 7156 61004 7162 61016
rect 7374 61004 7380 61016
rect 7432 61004 7438 61056
rect 8386 61004 8392 61056
rect 8444 61004 8450 61056
rect 1104 60954 8832 60976
rect 1104 60902 3010 60954
rect 3062 60902 3074 60954
rect 3126 60902 3138 60954
rect 3190 60902 3202 60954
rect 3254 60902 3266 60954
rect 3318 60902 8010 60954
rect 8062 60902 8074 60954
rect 8126 60902 8138 60954
rect 8190 60902 8202 60954
rect 8254 60902 8266 60954
rect 8318 60902 8832 60954
rect 1104 60880 8832 60902
rect 4706 60800 4712 60852
rect 4764 60840 4770 60852
rect 4801 60843 4859 60849
rect 4801 60840 4813 60843
rect 4764 60812 4813 60840
rect 4764 60800 4770 60812
rect 4801 60809 4813 60812
rect 4847 60809 4859 60843
rect 4801 60803 4859 60809
rect 5537 60843 5595 60849
rect 5537 60809 5549 60843
rect 5583 60840 5595 60843
rect 6086 60840 6092 60852
rect 5583 60812 6092 60840
rect 5583 60809 5595 60812
rect 5537 60803 5595 60809
rect 6086 60800 6092 60812
rect 6144 60800 6150 60852
rect 7098 60840 7104 60852
rect 6932 60812 7104 60840
rect 6932 60784 6960 60812
rect 7098 60800 7104 60812
rect 7156 60840 7162 60852
rect 7156 60812 7328 60840
rect 7156 60800 7162 60812
rect 6914 60732 6920 60784
rect 6972 60732 6978 60784
rect 7006 60732 7012 60784
rect 7064 60732 7070 60784
rect 7300 60772 7328 60812
rect 7374 60800 7380 60852
rect 7432 60840 7438 60852
rect 8018 60840 8024 60852
rect 7432 60812 8024 60840
rect 7432 60800 7438 60812
rect 8018 60800 8024 60812
rect 8076 60800 8082 60852
rect 7300 60744 7498 60772
rect 4985 60707 5043 60713
rect 4985 60673 4997 60707
rect 5031 60673 5043 60707
rect 4985 60667 5043 60673
rect 5000 60568 5028 60667
rect 5626 60664 5632 60716
rect 5684 60664 5690 60716
rect 5813 60639 5871 60645
rect 5813 60605 5825 60639
rect 5859 60636 5871 60639
rect 5902 60636 5908 60648
rect 5859 60608 5908 60636
rect 5859 60605 5871 60608
rect 5813 60599 5871 60605
rect 5902 60596 5908 60608
rect 5960 60596 5966 60648
rect 6730 60596 6736 60648
rect 6788 60596 6794 60648
rect 7006 60596 7012 60648
rect 7064 60636 7070 60648
rect 7374 60636 7380 60648
rect 7064 60608 7380 60636
rect 7064 60596 7070 60608
rect 7374 60596 7380 60608
rect 7432 60596 7438 60648
rect 5169 60571 5227 60577
rect 5169 60568 5181 60571
rect 5000 60540 5181 60568
rect 5169 60537 5181 60540
rect 5215 60537 5227 60571
rect 5169 60531 5227 60537
rect 7006 60460 7012 60512
rect 7064 60500 7070 60512
rect 7742 60500 7748 60512
rect 7064 60472 7748 60500
rect 7064 60460 7070 60472
rect 7742 60460 7748 60472
rect 7800 60500 7806 60512
rect 8481 60503 8539 60509
rect 8481 60500 8493 60503
rect 7800 60472 8493 60500
rect 7800 60460 7806 60472
rect 8481 60469 8493 60472
rect 8527 60469 8539 60503
rect 8481 60463 8539 60469
rect 1104 60410 8832 60432
rect 1104 60358 2350 60410
rect 2402 60358 2414 60410
rect 2466 60358 2478 60410
rect 2530 60358 2542 60410
rect 2594 60358 2606 60410
rect 2658 60358 7350 60410
rect 7402 60358 7414 60410
rect 7466 60358 7478 60410
rect 7530 60358 7542 60410
rect 7594 60358 7606 60410
rect 7658 60358 8832 60410
rect 1104 60336 8832 60358
rect 6641 60299 6699 60305
rect 6641 60265 6653 60299
rect 6687 60296 6699 60299
rect 6822 60296 6828 60308
rect 6687 60268 6828 60296
rect 6687 60265 6699 60268
rect 6641 60259 6699 60265
rect 6822 60256 6828 60268
rect 6880 60256 6886 60308
rect 5169 60231 5227 60237
rect 5169 60197 5181 60231
rect 5215 60197 5227 60231
rect 5169 60191 5227 60197
rect 5077 60095 5135 60101
rect 5077 60061 5089 60095
rect 5123 60092 5135 60095
rect 5184 60092 5212 60191
rect 5813 60163 5871 60169
rect 5813 60129 5825 60163
rect 5859 60160 5871 60163
rect 5902 60160 5908 60172
rect 5859 60132 5908 60160
rect 5859 60129 5871 60132
rect 5813 60123 5871 60129
rect 5902 60120 5908 60132
rect 5960 60120 5966 60172
rect 7193 60163 7251 60169
rect 7193 60129 7205 60163
rect 7239 60160 7251 60163
rect 8018 60160 8024 60172
rect 7239 60132 8024 60160
rect 7239 60129 7251 60132
rect 7193 60123 7251 60129
rect 5123 60064 5212 60092
rect 5123 60061 5135 60064
rect 5077 60055 5135 60061
rect 7006 60052 7012 60104
rect 7064 60052 7070 60104
rect 5537 60027 5595 60033
rect 5537 59993 5549 60027
rect 5583 60024 5595 60027
rect 5718 60024 5724 60036
rect 5583 59996 5724 60024
rect 5583 59993 5595 59996
rect 5537 59987 5595 59993
rect 5718 59984 5724 59996
rect 5776 60024 5782 60036
rect 7101 60027 7159 60033
rect 7101 60024 7113 60027
rect 5776 59996 7113 60024
rect 5776 59984 5782 59996
rect 7101 59993 7113 59996
rect 7147 59993 7159 60027
rect 7101 59987 7159 59993
rect 4890 59916 4896 59968
rect 4948 59916 4954 59968
rect 5629 59959 5687 59965
rect 5629 59925 5641 59959
rect 5675 59956 5687 59959
rect 6178 59956 6184 59968
rect 5675 59928 6184 59956
rect 5675 59925 5687 59928
rect 5629 59919 5687 59925
rect 6178 59916 6184 59928
rect 6236 59916 6242 59968
rect 7006 59916 7012 59968
rect 7064 59956 7070 59968
rect 7208 59956 7236 60123
rect 8018 60120 8024 60132
rect 8076 60120 8082 60172
rect 7742 60052 7748 60104
rect 7800 60092 7806 60104
rect 8205 60095 8263 60101
rect 8205 60092 8217 60095
rect 7800 60064 8217 60092
rect 7800 60052 7806 60064
rect 8205 60061 8217 60064
rect 8251 60061 8263 60095
rect 8205 60055 8263 60061
rect 7064 59928 7236 59956
rect 7064 59916 7070 59928
rect 8386 59916 8392 59968
rect 8444 59916 8450 59968
rect 1104 59866 8832 59888
rect 1104 59814 3010 59866
rect 3062 59814 3074 59866
rect 3126 59814 3138 59866
rect 3190 59814 3202 59866
rect 3254 59814 3266 59866
rect 3318 59814 8010 59866
rect 8062 59814 8074 59866
rect 8126 59814 8138 59866
rect 8190 59814 8202 59866
rect 8254 59814 8266 59866
rect 8318 59814 8832 59866
rect 1104 59792 8832 59814
rect 4890 59752 4896 59764
rect 4724 59724 4896 59752
rect 4724 59693 4752 59724
rect 4890 59712 4896 59724
rect 4948 59712 4954 59764
rect 6641 59755 6699 59761
rect 6641 59721 6653 59755
rect 6687 59721 6699 59755
rect 6641 59715 6699 59721
rect 4709 59687 4767 59693
rect 4709 59653 4721 59687
rect 4755 59653 4767 59687
rect 6656 59684 6684 59715
rect 7009 59687 7067 59693
rect 7009 59684 7021 59687
rect 6656 59656 7021 59684
rect 4709 59647 4767 59653
rect 7009 59653 7021 59656
rect 7055 59653 7067 59687
rect 7009 59647 7067 59653
rect 4430 59576 4436 59628
rect 4488 59576 4494 59628
rect 5736 59588 5842 59616
rect 5736 59480 5764 59588
rect 6454 59576 6460 59628
rect 6512 59576 6518 59628
rect 6730 59508 6736 59560
rect 6788 59508 6794 59560
rect 7098 59548 7104 59560
rect 6840 59520 7104 59548
rect 6840 59480 6868 59520
rect 7098 59508 7104 59520
rect 7156 59548 7162 59560
rect 8128 59548 8156 59602
rect 7156 59520 8156 59548
rect 7156 59508 7162 59520
rect 5736 59452 6868 59480
rect 5736 59424 5764 59452
rect 5718 59372 5724 59424
rect 5776 59372 5782 59424
rect 6178 59372 6184 59424
rect 6236 59372 6242 59424
rect 7098 59372 7104 59424
rect 7156 59412 7162 59424
rect 7742 59412 7748 59424
rect 7156 59384 7748 59412
rect 7156 59372 7162 59384
rect 7742 59372 7748 59384
rect 7800 59412 7806 59424
rect 8481 59415 8539 59421
rect 8481 59412 8493 59415
rect 7800 59384 8493 59412
rect 7800 59372 7806 59384
rect 8481 59381 8493 59384
rect 8527 59381 8539 59415
rect 8481 59375 8539 59381
rect 1104 59322 8832 59344
rect 1104 59270 2350 59322
rect 2402 59270 2414 59322
rect 2466 59270 2478 59322
rect 2530 59270 2542 59322
rect 2594 59270 2606 59322
rect 2658 59270 7350 59322
rect 7402 59270 7414 59322
rect 7466 59270 7478 59322
rect 7530 59270 7542 59322
rect 7594 59270 7606 59322
rect 7658 59270 8832 59322
rect 1104 59248 8832 59270
rect 6454 59168 6460 59220
rect 6512 59208 6518 59220
rect 6733 59211 6791 59217
rect 6733 59208 6745 59211
rect 6512 59180 6745 59208
rect 6512 59168 6518 59180
rect 6733 59177 6745 59180
rect 6779 59177 6791 59211
rect 6733 59171 6791 59177
rect 7006 59100 7012 59152
rect 7064 59140 7070 59152
rect 7064 59112 7420 59140
rect 7064 59100 7070 59112
rect 5902 59032 5908 59084
rect 5960 59032 5966 59084
rect 6178 59032 6184 59084
rect 6236 59072 6242 59084
rect 7392 59081 7420 59112
rect 7193 59075 7251 59081
rect 7193 59072 7205 59075
rect 6236 59044 7205 59072
rect 6236 59032 6242 59044
rect 7193 59041 7205 59044
rect 7239 59041 7251 59075
rect 7193 59035 7251 59041
rect 7377 59075 7435 59081
rect 7377 59041 7389 59075
rect 7423 59041 7435 59075
rect 7377 59035 7435 59041
rect 5629 59007 5687 59013
rect 5629 58973 5641 59007
rect 5675 59004 5687 59007
rect 6196 59004 6224 59032
rect 5675 58976 6224 59004
rect 5675 58973 5687 58976
rect 5629 58967 5687 58973
rect 7098 58964 7104 59016
rect 7156 58964 7162 59016
rect 7742 58896 7748 58948
rect 7800 58936 7806 58948
rect 8113 58939 8171 58945
rect 8113 58936 8125 58939
rect 7800 58908 8125 58936
rect 7800 58896 7806 58908
rect 8113 58905 8125 58908
rect 8159 58905 8171 58939
rect 8113 58899 8171 58905
rect 5258 58828 5264 58880
rect 5316 58828 5322 58880
rect 5721 58871 5779 58877
rect 5721 58837 5733 58871
rect 5767 58868 5779 58871
rect 5994 58868 6000 58880
rect 5767 58840 6000 58868
rect 5767 58837 5779 58840
rect 5721 58831 5779 58837
rect 5994 58828 6000 58840
rect 6052 58828 6058 58880
rect 8389 58871 8447 58877
rect 8389 58837 8401 58871
rect 8435 58868 8447 58871
rect 8478 58868 8484 58880
rect 8435 58840 8484 58868
rect 8435 58837 8447 58840
rect 8389 58831 8447 58837
rect 8478 58828 8484 58840
rect 8536 58828 8542 58880
rect 1104 58778 8832 58800
rect 1104 58726 3010 58778
rect 3062 58726 3074 58778
rect 3126 58726 3138 58778
rect 3190 58726 3202 58778
rect 3254 58726 3266 58778
rect 3318 58726 8010 58778
rect 8062 58726 8074 58778
rect 8126 58726 8138 58778
rect 8190 58726 8202 58778
rect 8254 58726 8266 58778
rect 8318 58726 8832 58778
rect 1104 58704 8832 58726
rect 5828 58636 7144 58664
rect 4706 58556 4712 58608
rect 4764 58556 4770 58608
rect 5718 58488 5724 58540
rect 5776 58528 5782 58540
rect 5828 58528 5856 58636
rect 7116 58596 7144 58636
rect 7116 58568 7498 58596
rect 5776 58514 5856 58528
rect 5776 58500 5842 58514
rect 5776 58488 5782 58500
rect 6454 58488 6460 58540
rect 6512 58488 6518 58540
rect 4433 58463 4491 58469
rect 4433 58429 4445 58463
rect 4479 58460 4491 58463
rect 6730 58460 6736 58472
rect 4479 58432 6736 58460
rect 4479 58429 4491 58432
rect 4433 58423 4491 58429
rect 6730 58420 6736 58432
rect 6788 58420 6794 58472
rect 7009 58463 7067 58469
rect 7009 58460 7021 58463
rect 6840 58432 7021 58460
rect 6641 58395 6699 58401
rect 6641 58361 6653 58395
rect 6687 58392 6699 58395
rect 6840 58392 6868 58432
rect 7009 58429 7021 58432
rect 7055 58429 7067 58463
rect 7009 58423 7067 58429
rect 6687 58364 6868 58392
rect 6687 58361 6699 58364
rect 6641 58355 6699 58361
rect 5994 58284 6000 58336
rect 6052 58324 6058 58336
rect 6181 58327 6239 58333
rect 6181 58324 6193 58327
rect 6052 58296 6193 58324
rect 6052 58284 6058 58296
rect 6181 58293 6193 58296
rect 6227 58293 6239 58327
rect 6181 58287 6239 58293
rect 7098 58284 7104 58336
rect 7156 58324 7162 58336
rect 7742 58324 7748 58336
rect 7156 58296 7748 58324
rect 7156 58284 7162 58296
rect 7742 58284 7748 58296
rect 7800 58324 7806 58336
rect 8481 58327 8539 58333
rect 8481 58324 8493 58327
rect 7800 58296 8493 58324
rect 7800 58284 7806 58296
rect 8481 58293 8493 58296
rect 8527 58293 8539 58327
rect 8481 58287 8539 58293
rect 1104 58234 8832 58256
rect 1104 58182 2350 58234
rect 2402 58182 2414 58234
rect 2466 58182 2478 58234
rect 2530 58182 2542 58234
rect 2594 58182 2606 58234
rect 2658 58182 7350 58234
rect 7402 58182 7414 58234
rect 7466 58182 7478 58234
rect 7530 58182 7542 58234
rect 7594 58182 7606 58234
rect 7658 58182 8832 58234
rect 1104 58160 8832 58182
rect 4706 58080 4712 58132
rect 4764 58120 4770 58132
rect 4985 58123 5043 58129
rect 4985 58120 4997 58123
rect 4764 58092 4997 58120
rect 4764 58080 4770 58092
rect 4985 58089 4997 58092
rect 5031 58089 5043 58123
rect 4985 58083 5043 58089
rect 6454 58080 6460 58132
rect 6512 58120 6518 58132
rect 6733 58123 6791 58129
rect 6733 58120 6745 58123
rect 6512 58092 6745 58120
rect 6512 58080 6518 58092
rect 6733 58089 6745 58092
rect 6779 58089 6791 58123
rect 6733 58083 6791 58089
rect 7006 57944 7012 57996
rect 7064 57984 7070 57996
rect 7377 57987 7435 57993
rect 7377 57984 7389 57987
rect 7064 57956 7389 57984
rect 7064 57944 7070 57956
rect 7377 57953 7389 57956
rect 7423 57984 7435 57987
rect 7742 57984 7748 57996
rect 7423 57956 7748 57984
rect 7423 57953 7435 57956
rect 7377 57947 7435 57953
rect 7742 57944 7748 57956
rect 7800 57944 7806 57996
rect 5169 57919 5227 57925
rect 5169 57885 5181 57919
rect 5215 57916 5227 57919
rect 5258 57916 5264 57928
rect 5215 57888 5264 57916
rect 5215 57885 5227 57888
rect 5169 57879 5227 57885
rect 5258 57876 5264 57888
rect 5316 57876 5322 57928
rect 7098 57876 7104 57928
rect 7156 57876 7162 57928
rect 6454 57808 6460 57860
rect 6512 57848 6518 57860
rect 8113 57851 8171 57857
rect 8113 57848 8125 57851
rect 6512 57820 8125 57848
rect 6512 57808 6518 57820
rect 8113 57817 8125 57820
rect 8159 57817 8171 57851
rect 8113 57811 8171 57817
rect 5994 57740 6000 57792
rect 6052 57780 6058 57792
rect 7193 57783 7251 57789
rect 7193 57780 7205 57783
rect 6052 57752 7205 57780
rect 6052 57740 6058 57752
rect 7193 57749 7205 57752
rect 7239 57749 7251 57783
rect 7193 57743 7251 57749
rect 7650 57740 7656 57792
rect 7708 57780 7714 57792
rect 8205 57783 8263 57789
rect 8205 57780 8217 57783
rect 7708 57752 8217 57780
rect 7708 57740 7714 57752
rect 8205 57749 8217 57752
rect 8251 57749 8263 57783
rect 8205 57743 8263 57749
rect 1104 57690 8832 57712
rect 1104 57638 3010 57690
rect 3062 57638 3074 57690
rect 3126 57638 3138 57690
rect 3190 57638 3202 57690
rect 3254 57638 3266 57690
rect 3318 57638 8010 57690
rect 8062 57638 8074 57690
rect 8126 57638 8138 57690
rect 8190 57638 8202 57690
rect 8254 57638 8266 57690
rect 8318 57638 8832 57690
rect 1104 57616 8832 57638
rect 5718 57468 5724 57520
rect 5776 57468 5782 57520
rect 6822 57400 6828 57452
rect 6880 57400 6886 57452
rect 7098 57400 7104 57452
rect 7156 57440 7162 57452
rect 7745 57443 7803 57449
rect 7745 57440 7757 57443
rect 7156 57412 7757 57440
rect 7156 57400 7162 57412
rect 7745 57409 7757 57412
rect 7791 57409 7803 57443
rect 7745 57403 7803 57409
rect 4433 57375 4491 57381
rect 4433 57341 4445 57375
rect 4479 57341 4491 57375
rect 4433 57335 4491 57341
rect 4448 57236 4476 57335
rect 4706 57332 4712 57384
rect 4764 57332 4770 57384
rect 7650 57332 7656 57384
rect 7708 57372 7714 57384
rect 8018 57372 8024 57384
rect 7708 57344 8024 57372
rect 7708 57332 7714 57344
rect 8018 57332 8024 57344
rect 8076 57332 8082 57384
rect 6086 57236 6092 57248
rect 4448 57208 6092 57236
rect 6086 57196 6092 57208
rect 6144 57196 6150 57248
rect 6178 57196 6184 57248
rect 6236 57196 6242 57248
rect 7006 57196 7012 57248
rect 7064 57196 7070 57248
rect 8021 57239 8079 57245
rect 8021 57205 8033 57239
rect 8067 57236 8079 57239
rect 8570 57236 8576 57248
rect 8067 57208 8576 57236
rect 8067 57205 8079 57208
rect 8021 57199 8079 57205
rect 8570 57196 8576 57208
rect 8628 57196 8634 57248
rect 1104 57146 8832 57168
rect 1104 57094 2350 57146
rect 2402 57094 2414 57146
rect 2466 57094 2478 57146
rect 2530 57094 2542 57146
rect 2594 57094 2606 57146
rect 2658 57094 7350 57146
rect 7402 57094 7414 57146
rect 7466 57094 7478 57146
rect 7530 57094 7542 57146
rect 7594 57094 7606 57146
rect 7658 57094 8832 57146
rect 1104 57072 8832 57094
rect 4706 56992 4712 57044
rect 4764 57032 4770 57044
rect 4801 57035 4859 57041
rect 4801 57032 4813 57035
rect 4764 57004 4813 57032
rect 4764 56992 4770 57004
rect 4801 57001 4813 57004
rect 4847 57001 4859 57035
rect 4801 56995 4859 57001
rect 5997 57035 6055 57041
rect 5997 57001 6009 57035
rect 6043 57032 6055 57035
rect 6270 57032 6276 57044
rect 6043 57004 6276 57032
rect 6043 57001 6055 57004
rect 5997 56995 6055 57001
rect 6270 56992 6276 57004
rect 6328 56992 6334 57044
rect 5077 56967 5135 56973
rect 5077 56933 5089 56967
rect 5123 56933 5135 56967
rect 6365 56967 6423 56973
rect 6365 56964 6377 56967
rect 5077 56927 5135 56933
rect 5920 56936 6377 56964
rect 4985 56831 5043 56837
rect 4985 56797 4997 56831
rect 5031 56828 5043 56831
rect 5092 56828 5120 56927
rect 5920 56908 5948 56936
rect 6365 56933 6377 56936
rect 6411 56933 6423 56967
rect 6365 56927 6423 56933
rect 5721 56899 5779 56905
rect 5721 56865 5733 56899
rect 5767 56896 5779 56899
rect 5902 56896 5908 56908
rect 5767 56868 5908 56896
rect 5767 56865 5779 56868
rect 5721 56859 5779 56865
rect 5902 56856 5908 56868
rect 5960 56856 5966 56908
rect 6086 56856 6092 56908
rect 6144 56896 6150 56908
rect 6730 56896 6736 56908
rect 6144 56868 6736 56896
rect 6144 56856 6150 56868
rect 6730 56856 6736 56868
rect 6788 56856 6794 56908
rect 7006 56856 7012 56908
rect 7064 56856 7070 56908
rect 7098 56856 7104 56908
rect 7156 56896 7162 56908
rect 8481 56899 8539 56905
rect 8481 56896 8493 56899
rect 7156 56868 8493 56896
rect 7156 56856 7162 56868
rect 8481 56865 8493 56868
rect 8527 56865 8539 56899
rect 8481 56859 8539 56865
rect 5031 56800 5120 56828
rect 5445 56831 5503 56837
rect 5031 56797 5043 56800
rect 4985 56791 5043 56797
rect 5445 56797 5457 56831
rect 5491 56828 5503 56831
rect 5994 56828 6000 56840
rect 5491 56800 6000 56828
rect 5491 56797 5503 56800
rect 5445 56791 5503 56797
rect 5994 56788 6000 56800
rect 6052 56788 6058 56840
rect 6181 56831 6239 56837
rect 6181 56797 6193 56831
rect 6227 56828 6239 56831
rect 6270 56828 6276 56840
rect 6227 56800 6276 56828
rect 6227 56797 6239 56800
rect 6181 56791 6239 56797
rect 6270 56788 6276 56800
rect 6328 56788 6334 56840
rect 8018 56788 8024 56840
rect 8076 56828 8082 56840
rect 8076 56814 8142 56828
rect 8076 56800 8156 56814
rect 8076 56788 8082 56800
rect 5537 56695 5595 56701
rect 5537 56661 5549 56695
rect 5583 56692 5595 56695
rect 5626 56692 5632 56704
rect 5583 56664 5632 56692
rect 5583 56661 5595 56664
rect 5537 56655 5595 56661
rect 5626 56652 5632 56664
rect 5684 56652 5690 56704
rect 7650 56652 7656 56704
rect 7708 56692 7714 56704
rect 8128 56692 8156 56800
rect 7708 56664 8156 56692
rect 7708 56652 7714 56664
rect 1104 56602 8832 56624
rect 1104 56550 3010 56602
rect 3062 56550 3074 56602
rect 3126 56550 3138 56602
rect 3190 56550 3202 56602
rect 3254 56550 3266 56602
rect 3318 56550 8010 56602
rect 8062 56550 8074 56602
rect 8126 56550 8138 56602
rect 8190 56550 8202 56602
rect 8254 56550 8266 56602
rect 8318 56550 8832 56602
rect 1104 56528 8832 56550
rect 5261 56491 5319 56497
rect 5261 56457 5273 56491
rect 5307 56457 5319 56491
rect 5261 56451 5319 56457
rect 5169 56355 5227 56361
rect 5169 56321 5181 56355
rect 5215 56352 5227 56355
rect 5276 56352 5304 56451
rect 6454 56448 6460 56500
rect 6512 56488 6518 56500
rect 6549 56491 6607 56497
rect 6549 56488 6561 56491
rect 6512 56460 6561 56488
rect 6512 56448 6518 56460
rect 6549 56457 6561 56460
rect 6595 56457 6607 56491
rect 6549 56451 6607 56457
rect 6733 56491 6791 56497
rect 6733 56457 6745 56491
rect 6779 56488 6791 56491
rect 6822 56488 6828 56500
rect 6779 56460 6828 56488
rect 6779 56457 6791 56460
rect 6733 56451 6791 56457
rect 6822 56448 6828 56460
rect 6880 56448 6886 56500
rect 7098 56448 7104 56500
rect 7156 56448 7162 56500
rect 5626 56380 5632 56432
rect 5684 56420 5690 56432
rect 6178 56420 6184 56432
rect 5684 56392 6184 56420
rect 5684 56380 5690 56392
rect 6178 56380 6184 56392
rect 6236 56420 6242 56432
rect 7193 56423 7251 56429
rect 7193 56420 7205 56423
rect 6236 56392 7205 56420
rect 6236 56380 6242 56392
rect 7193 56389 7205 56392
rect 7239 56389 7251 56423
rect 7193 56383 7251 56389
rect 5215 56324 5304 56352
rect 5215 56321 5227 56324
rect 5169 56315 5227 56321
rect 6362 56312 6368 56364
rect 6420 56352 6426 56364
rect 6457 56355 6515 56361
rect 6457 56352 6469 56355
rect 6420 56324 6469 56352
rect 6420 56312 6426 56324
rect 6457 56321 6469 56324
rect 6503 56321 6515 56355
rect 6457 56315 6515 56321
rect 5626 56244 5632 56296
rect 5684 56284 5690 56296
rect 5721 56287 5779 56293
rect 5721 56284 5733 56287
rect 5684 56256 5733 56284
rect 5684 56244 5690 56256
rect 5721 56253 5733 56256
rect 5767 56253 5779 56287
rect 5721 56247 5779 56253
rect 5902 56244 5908 56296
rect 5960 56244 5966 56296
rect 6914 56244 6920 56296
rect 6972 56284 6978 56296
rect 7285 56287 7343 56293
rect 7285 56284 7297 56287
rect 6972 56256 7297 56284
rect 6972 56244 6978 56256
rect 7285 56253 7297 56256
rect 7331 56284 7343 56287
rect 7742 56284 7748 56296
rect 7331 56256 7748 56284
rect 7331 56253 7343 56256
rect 7285 56247 7343 56253
rect 7742 56244 7748 56256
rect 7800 56244 7806 56296
rect 6822 56176 6828 56228
rect 6880 56216 6886 56228
rect 7926 56216 7932 56228
rect 6880 56188 7932 56216
rect 6880 56176 6886 56188
rect 7926 56176 7932 56188
rect 7984 56176 7990 56228
rect 4890 56108 4896 56160
rect 4948 56148 4954 56160
rect 4985 56151 5043 56157
rect 4985 56148 4997 56151
rect 4948 56120 4997 56148
rect 4948 56108 4954 56120
rect 4985 56117 4997 56120
rect 5031 56117 5043 56151
rect 4985 56111 5043 56117
rect 7650 56108 7656 56160
rect 7708 56148 7714 56160
rect 8018 56148 8024 56160
rect 7708 56120 8024 56148
rect 7708 56108 7714 56120
rect 8018 56108 8024 56120
rect 8076 56108 8082 56160
rect 1104 56058 8832 56080
rect 1104 56006 2350 56058
rect 2402 56006 2414 56058
rect 2466 56006 2478 56058
rect 2530 56006 2542 56058
rect 2594 56006 2606 56058
rect 2658 56006 7350 56058
rect 7402 56006 7414 56058
rect 7466 56006 7478 56058
rect 7530 56006 7542 56058
rect 7594 56006 7606 56058
rect 7658 56006 8832 56058
rect 1104 55984 8832 56006
rect 6454 55836 6460 55888
rect 6512 55836 6518 55888
rect 4801 55811 4859 55817
rect 4801 55777 4813 55811
rect 4847 55808 4859 55811
rect 4890 55808 4896 55820
rect 4847 55780 4896 55808
rect 4847 55777 4859 55780
rect 4801 55771 4859 55777
rect 4890 55768 4896 55780
rect 4948 55768 4954 55820
rect 6472 55808 6500 55836
rect 5920 55780 6500 55808
rect 5920 55752 5948 55780
rect 6730 55768 6736 55820
rect 6788 55768 6794 55820
rect 4430 55700 4436 55752
rect 4488 55740 4494 55752
rect 4525 55743 4583 55749
rect 4525 55740 4537 55743
rect 4488 55712 4537 55740
rect 4488 55700 4494 55712
rect 4525 55709 4537 55712
rect 4571 55709 4583 55743
rect 4525 55703 4583 55709
rect 5902 55700 5908 55752
rect 5960 55700 5966 55752
rect 6454 55700 6460 55752
rect 6512 55700 6518 55752
rect 8018 55700 8024 55752
rect 8076 55740 8082 55752
rect 8076 55712 8142 55740
rect 8076 55700 8082 55712
rect 7009 55675 7067 55681
rect 7009 55641 7021 55675
rect 7055 55641 7067 55675
rect 7009 55635 7067 55641
rect 5626 55564 5632 55616
rect 5684 55604 5690 55616
rect 6270 55604 6276 55616
rect 5684 55576 6276 55604
rect 5684 55564 5690 55576
rect 6270 55564 6276 55576
rect 6328 55564 6334 55616
rect 6641 55607 6699 55613
rect 6641 55573 6653 55607
rect 6687 55604 6699 55607
rect 7024 55604 7052 55635
rect 6687 55576 7052 55604
rect 6687 55573 6699 55576
rect 6641 55567 6699 55573
rect 8478 55564 8484 55616
rect 8536 55564 8542 55616
rect 1104 55514 8832 55536
rect 1104 55462 3010 55514
rect 3062 55462 3074 55514
rect 3126 55462 3138 55514
rect 3190 55462 3202 55514
rect 3254 55462 3266 55514
rect 3318 55462 8010 55514
rect 8062 55462 8074 55514
rect 8126 55462 8138 55514
rect 8190 55462 8202 55514
rect 8254 55462 8266 55514
rect 8318 55462 8832 55514
rect 1104 55440 8832 55462
rect 6270 55360 6276 55412
rect 6328 55360 6334 55412
rect 6454 55360 6460 55412
rect 6512 55400 6518 55412
rect 6641 55403 6699 55409
rect 6641 55400 6653 55403
rect 6512 55372 6653 55400
rect 6512 55360 6518 55372
rect 6641 55369 6653 55372
rect 6687 55369 6699 55403
rect 6641 55363 6699 55369
rect 6288 55332 6316 55360
rect 7101 55335 7159 55341
rect 7101 55332 7113 55335
rect 6288 55304 7113 55332
rect 7101 55301 7113 55304
rect 7147 55301 7159 55335
rect 7101 55295 7159 55301
rect 6270 55224 6276 55276
rect 6328 55264 6334 55276
rect 6638 55264 6644 55276
rect 6328 55236 6644 55264
rect 6328 55224 6334 55236
rect 6638 55224 6644 55236
rect 6696 55224 6702 55276
rect 7009 55267 7067 55273
rect 7009 55233 7021 55267
rect 7055 55264 7067 55267
rect 7837 55267 7895 55273
rect 7837 55264 7849 55267
rect 7055 55236 7849 55264
rect 7055 55233 7067 55236
rect 7009 55227 7067 55233
rect 7837 55233 7849 55236
rect 7883 55233 7895 55267
rect 7837 55227 7895 55233
rect 8478 55224 8484 55276
rect 8536 55224 8542 55276
rect 6914 55156 6920 55208
rect 6972 55196 6978 55208
rect 7193 55199 7251 55205
rect 7193 55196 7205 55199
rect 6972 55168 7205 55196
rect 6972 55156 6978 55168
rect 7193 55165 7205 55168
rect 7239 55165 7251 55199
rect 7193 55159 7251 55165
rect 1104 54970 8832 54992
rect 1104 54918 2350 54970
rect 2402 54918 2414 54970
rect 2466 54918 2478 54970
rect 2530 54918 2542 54970
rect 2594 54918 2606 54970
rect 2658 54918 7350 54970
rect 7402 54918 7414 54970
rect 7466 54918 7478 54970
rect 7530 54918 7542 54970
rect 7594 54918 7606 54970
rect 7658 54918 8832 54970
rect 1104 54896 8832 54918
rect 7561 54859 7619 54865
rect 7561 54825 7573 54859
rect 7607 54856 7619 54859
rect 8202 54856 8208 54868
rect 7607 54828 8208 54856
rect 7607 54825 7619 54828
rect 7561 54819 7619 54825
rect 8202 54816 8208 54828
rect 8260 54816 8266 54868
rect 7650 54748 7656 54800
rect 7708 54788 7714 54800
rect 7926 54788 7932 54800
rect 7708 54760 7932 54788
rect 7708 54748 7714 54760
rect 7926 54748 7932 54760
rect 7984 54748 7990 54800
rect 4430 54612 4436 54664
rect 4488 54652 4494 54664
rect 4525 54655 4583 54661
rect 4525 54652 4537 54655
rect 4488 54624 4537 54652
rect 4488 54612 4494 54624
rect 4525 54621 4537 54624
rect 4571 54621 4583 54655
rect 4525 54615 4583 54621
rect 5902 54612 5908 54664
rect 5960 54612 5966 54664
rect 7926 54612 7932 54664
rect 7984 54652 7990 54664
rect 8205 54655 8263 54661
rect 8205 54652 8217 54655
rect 7984 54624 8217 54652
rect 7984 54612 7990 54624
rect 8205 54621 8217 54624
rect 8251 54621 8263 54655
rect 8205 54615 8263 54621
rect 8478 54612 8484 54664
rect 8536 54612 8542 54664
rect 4798 54544 4804 54596
rect 4856 54544 4862 54596
rect 7653 54587 7711 54593
rect 7653 54553 7665 54587
rect 7699 54584 7711 54587
rect 8496 54584 8524 54612
rect 7699 54556 8524 54584
rect 7699 54553 7711 54556
rect 7653 54547 7711 54553
rect 5810 54476 5816 54528
rect 5868 54516 5874 54528
rect 6273 54519 6331 54525
rect 6273 54516 6285 54519
rect 5868 54488 6285 54516
rect 5868 54476 5874 54488
rect 6273 54485 6285 54488
rect 6319 54485 6331 54519
rect 6273 54479 6331 54485
rect 8386 54476 8392 54528
rect 8444 54476 8450 54528
rect 1104 54426 8832 54448
rect 1104 54374 3010 54426
rect 3062 54374 3074 54426
rect 3126 54374 3138 54426
rect 3190 54374 3202 54426
rect 3254 54374 3266 54426
rect 3318 54374 8010 54426
rect 8062 54374 8074 54426
rect 8126 54374 8138 54426
rect 8190 54374 8202 54426
rect 8254 54374 8266 54426
rect 8318 54374 8832 54426
rect 1104 54352 8832 54374
rect 4798 54272 4804 54324
rect 4856 54312 4862 54324
rect 4985 54315 5043 54321
rect 4985 54312 4997 54315
rect 4856 54284 4997 54312
rect 4856 54272 4862 54284
rect 4985 54281 4997 54284
rect 5031 54281 5043 54315
rect 4985 54275 5043 54281
rect 5261 54315 5319 54321
rect 5261 54281 5273 54315
rect 5307 54281 5319 54315
rect 5261 54275 5319 54281
rect 5169 54179 5227 54185
rect 5169 54145 5181 54179
rect 5215 54176 5227 54179
rect 5276 54176 5304 54275
rect 5626 54272 5632 54324
rect 5684 54272 5690 54324
rect 7650 54204 7656 54256
rect 7708 54204 7714 54256
rect 5215 54148 5304 54176
rect 5215 54145 5227 54148
rect 5169 54139 5227 54145
rect 6454 54136 6460 54188
rect 6512 54136 6518 54188
rect 6730 54136 6736 54188
rect 6788 54136 6794 54188
rect 5721 54111 5779 54117
rect 5721 54077 5733 54111
rect 5767 54077 5779 54111
rect 5721 54071 5779 54077
rect 5905 54111 5963 54117
rect 5905 54077 5917 54111
rect 5951 54108 5963 54111
rect 6178 54108 6184 54120
rect 5951 54080 6184 54108
rect 5951 54077 5963 54080
rect 5905 54071 5963 54077
rect 5736 53972 5764 54071
rect 6178 54068 6184 54080
rect 6236 54068 6242 54120
rect 7009 54111 7067 54117
rect 7009 54108 7021 54111
rect 6656 54080 7021 54108
rect 6656 54049 6684 54080
rect 7009 54077 7021 54080
rect 7055 54077 7067 54111
rect 7009 54071 7067 54077
rect 7650 54068 7656 54120
rect 7708 54108 7714 54120
rect 7708 54080 8064 54108
rect 7708 54068 7714 54080
rect 6641 54043 6699 54049
rect 6641 54009 6653 54043
rect 6687 54009 6699 54043
rect 8036 54040 8064 54080
rect 8110 54040 8116 54052
rect 8036 54012 8116 54040
rect 6641 54003 6699 54009
rect 8110 54000 8116 54012
rect 8168 54000 8174 54052
rect 5810 53972 5816 53984
rect 5736 53944 5816 53972
rect 5810 53932 5816 53944
rect 5868 53932 5874 53984
rect 7006 53932 7012 53984
rect 7064 53972 7070 53984
rect 8018 53972 8024 53984
rect 7064 53944 8024 53972
rect 7064 53932 7070 53944
rect 8018 53932 8024 53944
rect 8076 53972 8082 53984
rect 8481 53975 8539 53981
rect 8481 53972 8493 53975
rect 8076 53944 8493 53972
rect 8076 53932 8082 53944
rect 8481 53941 8493 53944
rect 8527 53941 8539 53975
rect 8481 53935 8539 53941
rect 1104 53882 8832 53904
rect 1104 53830 2350 53882
rect 2402 53830 2414 53882
rect 2466 53830 2478 53882
rect 2530 53830 2542 53882
rect 2594 53830 2606 53882
rect 2658 53830 7350 53882
rect 7402 53830 7414 53882
rect 7466 53830 7478 53882
rect 7530 53830 7542 53882
rect 7594 53830 7606 53882
rect 7658 53830 8832 53882
rect 1104 53808 8832 53830
rect 6454 53728 6460 53780
rect 6512 53768 6518 53780
rect 6641 53771 6699 53777
rect 6641 53768 6653 53771
rect 6512 53740 6653 53768
rect 6512 53728 6518 53740
rect 6641 53737 6653 53740
rect 6687 53737 6699 53771
rect 6641 53731 6699 53737
rect 5905 53635 5963 53641
rect 5905 53601 5917 53635
rect 5951 53632 5963 53635
rect 6178 53632 6184 53644
rect 5951 53604 6184 53632
rect 5951 53601 5963 53604
rect 5905 53595 5963 53601
rect 6178 53592 6184 53604
rect 6236 53632 6242 53644
rect 6638 53632 6644 53644
rect 6236 53604 6644 53632
rect 6236 53592 6242 53604
rect 6638 53592 6644 53604
rect 6696 53592 6702 53644
rect 6914 53592 6920 53644
rect 6972 53632 6978 53644
rect 7193 53635 7251 53641
rect 7193 53632 7205 53635
rect 6972 53604 7205 53632
rect 6972 53592 6978 53604
rect 7193 53601 7205 53604
rect 7239 53601 7251 53635
rect 7193 53595 7251 53601
rect 5169 53567 5227 53573
rect 5169 53533 5181 53567
rect 5215 53564 5227 53567
rect 5215 53536 5304 53564
rect 5215 53533 5227 53536
rect 5169 53527 5227 53533
rect 4982 53388 4988 53440
rect 5040 53388 5046 53440
rect 5276 53437 5304 53536
rect 7006 53524 7012 53576
rect 7064 53524 7070 53576
rect 5629 53499 5687 53505
rect 5629 53465 5641 53499
rect 5675 53496 5687 53499
rect 5810 53496 5816 53508
rect 5675 53468 5816 53496
rect 5675 53465 5687 53468
rect 5629 53459 5687 53465
rect 5810 53456 5816 53468
rect 5868 53496 5874 53508
rect 7101 53499 7159 53505
rect 7101 53496 7113 53499
rect 5868 53468 7113 53496
rect 5868 53456 5874 53468
rect 7101 53465 7113 53468
rect 7147 53465 7159 53499
rect 7101 53459 7159 53465
rect 5261 53431 5319 53437
rect 5261 53397 5273 53431
rect 5307 53397 5319 53431
rect 5261 53391 5319 53397
rect 5721 53431 5779 53437
rect 5721 53397 5733 53431
rect 5767 53428 5779 53431
rect 6178 53428 6184 53440
rect 5767 53400 6184 53428
rect 5767 53397 5779 53400
rect 5721 53391 5779 53397
rect 6178 53388 6184 53400
rect 6236 53388 6242 53440
rect 1104 53338 8832 53360
rect 1104 53286 3010 53338
rect 3062 53286 3074 53338
rect 3126 53286 3138 53338
rect 3190 53286 3202 53338
rect 3254 53286 3266 53338
rect 3318 53286 8010 53338
rect 8062 53286 8074 53338
rect 8126 53286 8138 53338
rect 8190 53286 8202 53338
rect 8254 53286 8266 53338
rect 8318 53286 8832 53338
rect 1104 53264 8832 53286
rect 4982 53224 4988 53236
rect 4724 53196 4988 53224
rect 4724 53165 4752 53196
rect 4982 53184 4988 53196
rect 5040 53184 5046 53236
rect 7926 53184 7932 53236
rect 7984 53224 7990 53236
rect 7984 53196 8156 53224
rect 7984 53184 7990 53196
rect 4709 53159 4767 53165
rect 4709 53125 4721 53159
rect 4755 53125 4767 53159
rect 4709 53119 4767 53125
rect 5842 53060 5948 53088
rect 5920 53032 5948 53060
rect 6454 53048 6460 53100
rect 6512 53048 6518 53100
rect 6730 53048 6736 53100
rect 6788 53048 6794 53100
rect 8128 53074 8156 53196
rect 4430 52980 4436 53032
rect 4488 52980 4494 53032
rect 5902 52980 5908 53032
rect 5960 52980 5966 53032
rect 7009 53023 7067 53029
rect 7009 53020 7021 53023
rect 6656 52992 7021 53020
rect 6656 52961 6684 52992
rect 7009 52989 7021 52992
rect 7055 52989 7067 53023
rect 7009 52983 7067 52989
rect 6641 52955 6699 52961
rect 6641 52921 6653 52955
rect 6687 52921 6699 52955
rect 6641 52915 6699 52921
rect 6178 52844 6184 52896
rect 6236 52844 6242 52896
rect 8202 52844 8208 52896
rect 8260 52884 8266 52896
rect 8481 52887 8539 52893
rect 8481 52884 8493 52887
rect 8260 52856 8493 52884
rect 8260 52844 8266 52856
rect 8481 52853 8493 52856
rect 8527 52853 8539 52887
rect 8481 52847 8539 52853
rect 1104 52794 8832 52816
rect 1104 52742 2350 52794
rect 2402 52742 2414 52794
rect 2466 52742 2478 52794
rect 2530 52742 2542 52794
rect 2594 52742 2606 52794
rect 2658 52742 7350 52794
rect 7402 52742 7414 52794
rect 7466 52742 7478 52794
rect 7530 52742 7542 52794
rect 7594 52742 7606 52794
rect 7658 52742 8832 52794
rect 1104 52720 8832 52742
rect 6454 52640 6460 52692
rect 6512 52680 6518 52692
rect 6641 52683 6699 52689
rect 6641 52680 6653 52683
rect 6512 52652 6653 52680
rect 6512 52640 6518 52652
rect 6641 52649 6653 52652
rect 6687 52649 6699 52683
rect 6641 52643 6699 52649
rect 8386 52640 8392 52692
rect 8444 52640 8450 52692
rect 6914 52572 6920 52624
rect 6972 52612 6978 52624
rect 6972 52584 7236 52612
rect 6972 52572 6978 52584
rect 7208 52553 7236 52584
rect 7101 52547 7159 52553
rect 7101 52544 7113 52547
rect 6196 52516 7113 52544
rect 6196 52488 6224 52516
rect 7101 52513 7113 52516
rect 7147 52513 7159 52547
rect 7101 52507 7159 52513
rect 7193 52547 7251 52553
rect 7193 52513 7205 52547
rect 7239 52513 7251 52547
rect 7193 52507 7251 52513
rect 6178 52436 6184 52488
rect 6236 52436 6242 52488
rect 7009 52479 7067 52485
rect 7009 52445 7021 52479
rect 7055 52476 7067 52479
rect 8202 52476 8208 52488
rect 7055 52448 8208 52476
rect 7055 52445 7067 52448
rect 7009 52439 7067 52445
rect 8202 52436 8208 52448
rect 8260 52436 8266 52488
rect 1104 52250 8832 52272
rect 1104 52198 3010 52250
rect 3062 52198 3074 52250
rect 3126 52198 3138 52250
rect 3190 52198 3202 52250
rect 3254 52198 3266 52250
rect 3318 52198 8010 52250
rect 8062 52198 8074 52250
rect 8126 52198 8138 52250
rect 8190 52198 8202 52250
rect 8254 52198 8266 52250
rect 8318 52198 8832 52250
rect 1104 52176 8832 52198
rect 7926 52096 7932 52148
rect 7984 52136 7990 52148
rect 8110 52136 8116 52148
rect 7984 52108 8116 52136
rect 7984 52096 7990 52108
rect 8110 52096 8116 52108
rect 8168 52096 8174 52148
rect 7944 52068 7972 52096
rect 5934 52040 7972 52068
rect 7926 51960 7932 52012
rect 7984 52000 7990 52012
rect 8205 52003 8263 52009
rect 8205 52000 8217 52003
rect 7984 51972 8217 52000
rect 7984 51960 7990 51972
rect 8205 51969 8217 51972
rect 8251 51969 8263 52003
rect 8205 51963 8263 51969
rect 4430 51892 4436 51944
rect 4488 51892 4494 51944
rect 4706 51892 4712 51944
rect 4764 51892 4770 51944
rect 5718 51756 5724 51808
rect 5776 51796 5782 51808
rect 6181 51799 6239 51805
rect 6181 51796 6193 51799
rect 5776 51768 6193 51796
rect 5776 51756 5782 51768
rect 6181 51765 6193 51768
rect 6227 51765 6239 51799
rect 6181 51759 6239 51765
rect 8386 51756 8392 51808
rect 8444 51756 8450 51808
rect 1104 51706 8832 51728
rect 1104 51654 2350 51706
rect 2402 51654 2414 51706
rect 2466 51654 2478 51706
rect 2530 51654 2542 51706
rect 2594 51654 2606 51706
rect 2658 51654 7350 51706
rect 7402 51654 7414 51706
rect 7466 51654 7478 51706
rect 7530 51654 7542 51706
rect 7594 51654 7606 51706
rect 7658 51654 8832 51706
rect 1104 51632 8832 51654
rect 4706 51552 4712 51604
rect 4764 51592 4770 51604
rect 4893 51595 4951 51601
rect 4893 51592 4905 51595
rect 4764 51564 4905 51592
rect 4764 51552 4770 51564
rect 4893 51561 4905 51564
rect 4939 51561 4951 51595
rect 4893 51555 4951 51561
rect 7098 51552 7104 51604
rect 7156 51592 7162 51604
rect 7374 51592 7380 51604
rect 7156 51564 7380 51592
rect 7156 51552 7162 51564
rect 7374 51552 7380 51564
rect 7432 51552 7438 51604
rect 5718 51416 5724 51468
rect 5776 51416 5782 51468
rect 5902 51416 5908 51468
rect 5960 51416 5966 51468
rect 6730 51416 6736 51468
rect 6788 51416 6794 51468
rect 7006 51416 7012 51468
rect 7064 51456 7070 51468
rect 7064 51428 8156 51456
rect 7064 51416 7070 51428
rect 8128 51400 8156 51428
rect 5077 51391 5135 51397
rect 5077 51357 5089 51391
rect 5123 51388 5135 51391
rect 5629 51391 5687 51397
rect 5123 51360 5304 51388
rect 5123 51357 5135 51360
rect 5077 51351 5135 51357
rect 5276 51261 5304 51360
rect 5629 51357 5641 51391
rect 5675 51388 5687 51391
rect 6178 51388 6184 51400
rect 5675 51360 6184 51388
rect 5675 51357 5687 51360
rect 5629 51351 5687 51357
rect 6178 51348 6184 51360
rect 6236 51348 6242 51400
rect 6454 51348 6460 51400
rect 6512 51348 6518 51400
rect 8110 51348 8116 51400
rect 8168 51348 8174 51400
rect 7009 51323 7067 51329
rect 7009 51289 7021 51323
rect 7055 51289 7067 51323
rect 7009 51283 7067 51289
rect 5261 51255 5319 51261
rect 5261 51221 5273 51255
rect 5307 51221 5319 51255
rect 5261 51215 5319 51221
rect 6641 51255 6699 51261
rect 6641 51221 6653 51255
rect 6687 51252 6699 51255
rect 7024 51252 7052 51283
rect 6687 51224 7052 51252
rect 6687 51221 6699 51224
rect 6641 51215 6699 51221
rect 7926 51212 7932 51264
rect 7984 51252 7990 51264
rect 8481 51255 8539 51261
rect 8481 51252 8493 51255
rect 7984 51224 8493 51252
rect 7984 51212 7990 51224
rect 8481 51221 8493 51224
rect 8527 51221 8539 51255
rect 8481 51215 8539 51221
rect 1104 51162 8832 51184
rect 1104 51110 3010 51162
rect 3062 51110 3074 51162
rect 3126 51110 3138 51162
rect 3190 51110 3202 51162
rect 3254 51110 3266 51162
rect 3318 51110 8010 51162
rect 8062 51110 8074 51162
rect 8126 51110 8138 51162
rect 8190 51110 8202 51162
rect 8254 51110 8266 51162
rect 8318 51110 8832 51162
rect 1104 51088 8832 51110
rect 5353 51051 5411 51057
rect 5353 51017 5365 51051
rect 5399 51017 5411 51051
rect 5353 51011 5411 51017
rect 5169 50915 5227 50921
rect 5169 50881 5181 50915
rect 5215 50912 5227 50915
rect 5368 50912 5396 51011
rect 6454 51008 6460 51060
rect 6512 51048 6518 51060
rect 6641 51051 6699 51057
rect 6641 51048 6653 51051
rect 6512 51020 6653 51048
rect 6512 51008 6518 51020
rect 6641 51017 6653 51020
rect 6687 51017 6699 51051
rect 6641 51011 6699 51017
rect 7009 51051 7067 51057
rect 7009 51017 7021 51051
rect 7055 51048 7067 51051
rect 7926 51048 7932 51060
rect 7055 51020 7932 51048
rect 7055 51017 7067 51020
rect 7009 51011 7067 51017
rect 7926 51008 7932 51020
rect 7984 51008 7990 51060
rect 5215 50884 5396 50912
rect 5215 50881 5227 50884
rect 5169 50875 5227 50881
rect 5718 50872 5724 50924
rect 5776 50912 5782 50924
rect 7101 50915 7159 50921
rect 7101 50912 7113 50915
rect 5776 50884 7113 50912
rect 5776 50872 5782 50884
rect 7101 50881 7113 50884
rect 7147 50881 7159 50915
rect 7101 50875 7159 50881
rect 5810 50804 5816 50856
rect 5868 50804 5874 50856
rect 5902 50804 5908 50856
rect 5960 50804 5966 50856
rect 6914 50804 6920 50856
rect 6972 50844 6978 50856
rect 7193 50847 7251 50853
rect 7193 50844 7205 50847
rect 6972 50816 7205 50844
rect 6972 50804 6978 50816
rect 7116 50720 7144 50816
rect 7193 50813 7205 50816
rect 7239 50813 7251 50847
rect 7193 50807 7251 50813
rect 4890 50668 4896 50720
rect 4948 50708 4954 50720
rect 4985 50711 5043 50717
rect 4985 50708 4997 50711
rect 4948 50680 4997 50708
rect 4948 50668 4954 50680
rect 4985 50677 4997 50680
rect 5031 50677 5043 50711
rect 4985 50671 5043 50677
rect 5718 50668 5724 50720
rect 5776 50708 5782 50720
rect 6546 50708 6552 50720
rect 5776 50680 6552 50708
rect 5776 50668 5782 50680
rect 6546 50668 6552 50680
rect 6604 50668 6610 50720
rect 7098 50668 7104 50720
rect 7156 50668 7162 50720
rect 7374 50668 7380 50720
rect 7432 50708 7438 50720
rect 7834 50708 7840 50720
rect 7432 50680 7840 50708
rect 7432 50668 7438 50680
rect 7834 50668 7840 50680
rect 7892 50668 7898 50720
rect 1104 50618 8832 50640
rect 1104 50566 2350 50618
rect 2402 50566 2414 50618
rect 2466 50566 2478 50618
rect 2530 50566 2542 50618
rect 2594 50566 2606 50618
rect 2658 50566 7350 50618
rect 7402 50566 7414 50618
rect 7466 50566 7478 50618
rect 7530 50566 7542 50618
rect 7594 50566 7606 50618
rect 7658 50566 8832 50618
rect 1104 50544 8832 50566
rect 5810 50464 5816 50516
rect 5868 50504 5874 50516
rect 6273 50507 6331 50513
rect 6273 50504 6285 50507
rect 5868 50476 6285 50504
rect 5868 50464 5874 50476
rect 6273 50473 6285 50476
rect 6319 50473 6331 50507
rect 6273 50467 6331 50473
rect 6641 50439 6699 50445
rect 6641 50405 6653 50439
rect 6687 50405 6699 50439
rect 6641 50399 6699 50405
rect 4801 50371 4859 50377
rect 4801 50337 4813 50371
rect 4847 50368 4859 50371
rect 4890 50368 4896 50380
rect 4847 50340 4896 50368
rect 4847 50337 4859 50340
rect 4801 50331 4859 50337
rect 4890 50328 4896 50340
rect 4948 50328 4954 50380
rect 6656 50368 6684 50399
rect 7009 50371 7067 50377
rect 7009 50368 7021 50371
rect 6656 50340 7021 50368
rect 7009 50337 7021 50340
rect 7055 50337 7067 50371
rect 7009 50331 7067 50337
rect 4430 50260 4436 50312
rect 4488 50300 4494 50312
rect 4525 50303 4583 50309
rect 4525 50300 4537 50303
rect 4488 50272 4537 50300
rect 4488 50260 4494 50272
rect 4525 50269 4537 50272
rect 4571 50269 4583 50303
rect 4525 50263 4583 50269
rect 6454 50260 6460 50312
rect 6512 50260 6518 50312
rect 6546 50260 6552 50312
rect 6604 50300 6610 50312
rect 6730 50300 6736 50312
rect 6604 50272 6736 50300
rect 6604 50260 6610 50272
rect 6730 50260 6736 50272
rect 6788 50260 6794 50312
rect 6026 50204 6592 50232
rect 6564 50164 6592 50204
rect 6914 50164 6920 50176
rect 6564 50136 6920 50164
rect 6914 50124 6920 50136
rect 6972 50164 6978 50176
rect 7926 50164 7932 50176
rect 6972 50136 7932 50164
rect 6972 50124 6978 50136
rect 7926 50124 7932 50136
rect 7984 50164 7990 50176
rect 8128 50164 8156 50286
rect 7984 50136 8156 50164
rect 8481 50167 8539 50173
rect 7984 50124 7990 50136
rect 8481 50133 8493 50167
rect 8527 50164 8539 50167
rect 8527 50136 8892 50164
rect 8527 50133 8539 50136
rect 8481 50127 8539 50133
rect 1104 50074 8832 50096
rect 1104 50022 3010 50074
rect 3062 50022 3074 50074
rect 3126 50022 3138 50074
rect 3190 50022 3202 50074
rect 3254 50022 3266 50074
rect 3318 50022 8010 50074
rect 8062 50022 8074 50074
rect 8126 50022 8138 50074
rect 8190 50022 8202 50074
rect 8254 50022 8266 50074
rect 8318 50022 8832 50074
rect 1104 50000 8832 50022
rect 8386 49920 8392 49972
rect 8444 49920 8450 49972
rect 5445 49827 5503 49833
rect 5445 49793 5457 49827
rect 5491 49824 5503 49827
rect 5534 49824 5540 49836
rect 5491 49796 5540 49824
rect 5491 49793 5503 49796
rect 5445 49787 5503 49793
rect 5534 49784 5540 49796
rect 5592 49824 5598 49836
rect 7469 49827 7527 49833
rect 7469 49824 7481 49827
rect 5592 49796 7481 49824
rect 5592 49784 5598 49796
rect 7469 49793 7481 49796
rect 7515 49793 7527 49827
rect 7469 49787 7527 49793
rect 8205 49827 8263 49833
rect 8205 49793 8217 49827
rect 8251 49824 8263 49827
rect 8864 49824 8892 50136
rect 8251 49796 8892 49824
rect 8251 49793 8263 49796
rect 8205 49787 8263 49793
rect 4430 49716 4436 49768
rect 4488 49756 4494 49768
rect 4617 49759 4675 49765
rect 4617 49756 4629 49759
rect 4488 49728 4629 49756
rect 4488 49716 4494 49728
rect 4617 49725 4629 49728
rect 4663 49725 4675 49759
rect 4617 49719 4675 49725
rect 6546 49716 6552 49768
rect 6604 49756 6610 49768
rect 6641 49759 6699 49765
rect 6641 49756 6653 49759
rect 6604 49728 6653 49756
rect 6604 49716 6610 49728
rect 6641 49725 6653 49728
rect 6687 49725 6699 49759
rect 8220 49756 8248 49787
rect 6641 49719 6699 49725
rect 7024 49728 8248 49756
rect 7024 49700 7052 49728
rect 7006 49648 7012 49700
rect 7064 49648 7070 49700
rect 1104 49530 8832 49552
rect 1104 49478 2350 49530
rect 2402 49478 2414 49530
rect 2466 49478 2478 49530
rect 2530 49478 2542 49530
rect 2594 49478 2606 49530
rect 2658 49478 7350 49530
rect 7402 49478 7414 49530
rect 7466 49478 7478 49530
rect 7530 49478 7542 49530
rect 7594 49478 7606 49530
rect 7658 49478 8832 49530
rect 1104 49456 8832 49478
rect 6454 49376 6460 49428
rect 6512 49416 6518 49428
rect 6641 49419 6699 49425
rect 6641 49416 6653 49419
rect 6512 49388 6653 49416
rect 6512 49376 6518 49388
rect 6641 49385 6653 49388
rect 6687 49385 6699 49419
rect 6641 49379 6699 49385
rect 7466 49376 7472 49428
rect 7524 49416 7530 49428
rect 7926 49416 7932 49428
rect 7524 49388 7932 49416
rect 7524 49376 7530 49388
rect 7926 49376 7932 49388
rect 7984 49376 7990 49428
rect 7484 49348 7512 49376
rect 6104 49320 7512 49348
rect 4430 49172 4436 49224
rect 4488 49212 4494 49224
rect 4709 49215 4767 49221
rect 4709 49212 4721 49215
rect 4488 49184 4721 49212
rect 4488 49172 4494 49184
rect 4709 49181 4721 49184
rect 4755 49181 4767 49215
rect 6104 49198 6132 49320
rect 7098 49240 7104 49292
rect 7156 49280 7162 49292
rect 7193 49283 7251 49289
rect 7193 49280 7205 49283
rect 7156 49252 7205 49280
rect 7156 49240 7162 49252
rect 7193 49249 7205 49252
rect 7239 49249 7251 49283
rect 7193 49243 7251 49249
rect 4709 49175 4767 49181
rect 7006 49172 7012 49224
rect 7064 49172 7070 49224
rect 7653 49215 7711 49221
rect 7653 49181 7665 49215
rect 7699 49212 7711 49215
rect 7742 49212 7748 49224
rect 7699 49184 7748 49212
rect 7699 49181 7711 49184
rect 7653 49175 7711 49181
rect 7742 49172 7748 49184
rect 7800 49172 7806 49224
rect 7926 49172 7932 49224
rect 7984 49212 7990 49224
rect 8205 49215 8263 49221
rect 8205 49212 8217 49215
rect 7984 49184 8217 49212
rect 7984 49172 7990 49184
rect 8205 49181 8217 49184
rect 8251 49181 8263 49215
rect 8205 49175 8263 49181
rect 4982 49104 4988 49156
rect 5040 49104 5046 49156
rect 5902 49036 5908 49088
rect 5960 49076 5966 49088
rect 6457 49079 6515 49085
rect 6457 49076 6469 49079
rect 5960 49048 6469 49076
rect 5960 49036 5966 49048
rect 6457 49045 6469 49048
rect 6503 49045 6515 49079
rect 6457 49039 6515 49045
rect 6638 49036 6644 49088
rect 6696 49076 6702 49088
rect 7101 49079 7159 49085
rect 7101 49076 7113 49079
rect 6696 49048 7113 49076
rect 6696 49036 6702 49048
rect 7101 49045 7113 49048
rect 7147 49045 7159 49079
rect 7101 49039 7159 49045
rect 7282 49036 7288 49088
rect 7340 49076 7346 49088
rect 7469 49079 7527 49085
rect 7469 49076 7481 49079
rect 7340 49048 7481 49076
rect 7340 49036 7346 49048
rect 7469 49045 7481 49048
rect 7515 49045 7527 49079
rect 7469 49039 7527 49045
rect 8386 49036 8392 49088
rect 8444 49036 8450 49088
rect 1104 48986 8832 49008
rect 1104 48934 3010 48986
rect 3062 48934 3074 48986
rect 3126 48934 3138 48986
rect 3190 48934 3202 48986
rect 3254 48934 3266 48986
rect 3318 48934 8010 48986
rect 8062 48934 8074 48986
rect 8126 48934 8138 48986
rect 8190 48934 8202 48986
rect 8254 48934 8266 48986
rect 8318 48934 8832 48986
rect 1104 48912 8832 48934
rect 4982 48832 4988 48884
rect 5040 48872 5046 48884
rect 5077 48875 5135 48881
rect 5077 48872 5089 48875
rect 5040 48844 5089 48872
rect 5040 48832 5046 48844
rect 5077 48841 5089 48844
rect 5123 48841 5135 48875
rect 5077 48835 5135 48841
rect 5445 48875 5503 48881
rect 5445 48841 5457 48875
rect 5491 48841 5503 48875
rect 5445 48835 5503 48841
rect 5261 48739 5319 48745
rect 5261 48705 5273 48739
rect 5307 48736 5319 48739
rect 5460 48736 5488 48835
rect 5810 48832 5816 48884
rect 5868 48872 5874 48884
rect 6638 48872 6644 48884
rect 5868 48844 6644 48872
rect 5868 48832 5874 48844
rect 6638 48832 6644 48844
rect 6696 48832 6702 48884
rect 7282 48872 7288 48884
rect 7024 48844 7288 48872
rect 7024 48813 7052 48844
rect 7282 48832 7288 48844
rect 7340 48832 7346 48884
rect 7009 48807 7067 48813
rect 7009 48773 7021 48807
rect 7055 48773 7067 48807
rect 7009 48767 7067 48773
rect 7466 48764 7472 48816
rect 7524 48764 7530 48816
rect 5307 48708 5488 48736
rect 5307 48705 5319 48708
rect 5261 48699 5319 48705
rect 5902 48628 5908 48680
rect 5960 48628 5966 48680
rect 5994 48628 6000 48680
rect 6052 48628 6058 48680
rect 6546 48628 6552 48680
rect 6604 48668 6610 48680
rect 6733 48671 6791 48677
rect 6733 48668 6745 48671
rect 6604 48640 6745 48668
rect 6604 48628 6610 48640
rect 6733 48637 6745 48640
rect 6779 48637 6791 48671
rect 6733 48631 6791 48637
rect 7098 48628 7104 48680
rect 7156 48668 7162 48680
rect 7650 48668 7656 48680
rect 7156 48640 7656 48668
rect 7156 48628 7162 48640
rect 7650 48628 7656 48640
rect 7708 48628 7714 48680
rect 8018 48492 8024 48544
rect 8076 48532 8082 48544
rect 8481 48535 8539 48541
rect 8481 48532 8493 48535
rect 8076 48504 8493 48532
rect 8076 48492 8082 48504
rect 8481 48501 8493 48504
rect 8527 48501 8539 48535
rect 8481 48495 8539 48501
rect 1104 48442 8832 48464
rect 1104 48390 2350 48442
rect 2402 48390 2414 48442
rect 2466 48390 2478 48442
rect 2530 48390 2542 48442
rect 2594 48390 2606 48442
rect 2658 48390 7350 48442
rect 7402 48390 7414 48442
rect 7466 48390 7478 48442
rect 7530 48390 7542 48442
rect 7594 48390 7606 48442
rect 7658 48390 8832 48442
rect 1104 48368 8832 48390
rect 7561 48331 7619 48337
rect 7561 48297 7573 48331
rect 7607 48328 7619 48331
rect 7742 48328 7748 48340
rect 7607 48300 7748 48328
rect 7607 48297 7619 48300
rect 7561 48291 7619 48297
rect 7742 48288 7748 48300
rect 7800 48288 7806 48340
rect 5445 48263 5503 48269
rect 5445 48229 5457 48263
rect 5491 48229 5503 48263
rect 5445 48223 5503 48229
rect 5353 48127 5411 48133
rect 5353 48093 5365 48127
rect 5399 48124 5411 48127
rect 5460 48124 5488 48223
rect 7098 48220 7104 48272
rect 7156 48220 7162 48272
rect 5994 48152 6000 48204
rect 6052 48152 6058 48204
rect 7009 48195 7067 48201
rect 7009 48161 7021 48195
rect 7055 48192 7067 48195
rect 7116 48192 7144 48220
rect 7055 48164 7144 48192
rect 7055 48161 7067 48164
rect 7009 48155 7067 48161
rect 5399 48096 5488 48124
rect 5813 48127 5871 48133
rect 5399 48093 5411 48096
rect 5353 48087 5411 48093
rect 5813 48093 5825 48127
rect 5859 48124 5871 48127
rect 5902 48124 5908 48136
rect 5859 48096 5908 48124
rect 5859 48093 5871 48096
rect 5813 48087 5871 48093
rect 5902 48084 5908 48096
rect 5960 48124 5966 48136
rect 7101 48127 7159 48133
rect 7101 48124 7113 48127
rect 5960 48096 7113 48124
rect 5960 48084 5966 48096
rect 7101 48093 7113 48096
rect 7147 48093 7159 48127
rect 7101 48087 7159 48093
rect 7193 48127 7251 48133
rect 7193 48093 7205 48127
rect 7239 48124 7251 48127
rect 8018 48124 8024 48136
rect 7239 48096 8024 48124
rect 7239 48093 7251 48096
rect 7193 48087 7251 48093
rect 8018 48084 8024 48096
rect 8076 48084 8082 48136
rect 4890 47948 4896 48000
rect 4948 47988 4954 48000
rect 5169 47991 5227 47997
rect 5169 47988 5181 47991
rect 4948 47960 5181 47988
rect 4948 47948 4954 47960
rect 5169 47957 5181 47960
rect 5215 47957 5227 47991
rect 5169 47951 5227 47957
rect 5905 47991 5963 47997
rect 5905 47957 5917 47991
rect 5951 47988 5963 47991
rect 6178 47988 6184 48000
rect 5951 47960 6184 47988
rect 5951 47957 5963 47960
rect 5905 47951 5963 47957
rect 6178 47948 6184 47960
rect 6236 47948 6242 48000
rect 1104 47898 8832 47920
rect 1104 47846 3010 47898
rect 3062 47846 3074 47898
rect 3126 47846 3138 47898
rect 3190 47846 3202 47898
rect 3254 47846 3266 47898
rect 3318 47846 8010 47898
rect 8062 47846 8074 47898
rect 8126 47846 8138 47898
rect 8190 47846 8202 47898
rect 8254 47846 8266 47898
rect 8318 47846 8832 47898
rect 1104 47824 8832 47846
rect 4890 47784 4896 47796
rect 4724 47756 4896 47784
rect 4724 47725 4752 47756
rect 4890 47744 4896 47756
rect 4948 47744 4954 47796
rect 6641 47787 6699 47793
rect 6641 47753 6653 47787
rect 6687 47753 6699 47787
rect 6641 47747 6699 47753
rect 4709 47719 4767 47725
rect 4709 47685 4721 47719
rect 4755 47685 4767 47719
rect 6086 47716 6092 47728
rect 5934 47688 6092 47716
rect 4709 47679 4767 47685
rect 6086 47676 6092 47688
rect 6144 47676 6150 47728
rect 6656 47716 6684 47747
rect 7009 47719 7067 47725
rect 7009 47716 7021 47719
rect 6656 47688 7021 47716
rect 7009 47685 7021 47688
rect 7055 47685 7067 47719
rect 7009 47679 7067 47685
rect 7098 47676 7104 47728
rect 7156 47716 7162 47728
rect 7156 47688 7498 47716
rect 7156 47676 7162 47688
rect 6454 47608 6460 47660
rect 6512 47608 6518 47660
rect 4430 47540 4436 47592
rect 4488 47540 4494 47592
rect 6546 47540 6552 47592
rect 6604 47580 6610 47592
rect 6733 47583 6791 47589
rect 6733 47580 6745 47583
rect 6604 47552 6745 47580
rect 6604 47540 6610 47552
rect 6733 47549 6745 47552
rect 6779 47549 6791 47583
rect 6733 47543 6791 47549
rect 6178 47404 6184 47456
rect 6236 47404 6242 47456
rect 8481 47447 8539 47453
rect 8481 47413 8493 47447
rect 8527 47444 8539 47447
rect 8527 47416 8892 47444
rect 8527 47413 8539 47416
rect 8481 47407 8539 47413
rect 1104 47354 8832 47376
rect 1104 47302 2350 47354
rect 2402 47302 2414 47354
rect 2466 47302 2478 47354
rect 2530 47302 2542 47354
rect 2594 47302 2606 47354
rect 2658 47302 7350 47354
rect 7402 47302 7414 47354
rect 7466 47302 7478 47354
rect 7530 47302 7542 47354
rect 7594 47302 7606 47354
rect 7658 47302 8832 47354
rect 1104 47280 8832 47302
rect 6454 47200 6460 47252
rect 6512 47240 6518 47252
rect 6825 47243 6883 47249
rect 6825 47240 6837 47243
rect 6512 47212 6837 47240
rect 6512 47200 6518 47212
rect 6825 47209 6837 47212
rect 6871 47209 6883 47243
rect 6825 47203 6883 47209
rect 7006 47200 7012 47252
rect 7064 47200 7070 47252
rect 8386 47200 8392 47252
rect 8444 47200 8450 47252
rect 7024 47172 7052 47200
rect 7024 47144 7420 47172
rect 7392 47116 7420 47144
rect 5994 47064 6000 47116
rect 6052 47064 6058 47116
rect 6178 47104 6184 47116
rect 6104 47076 6184 47104
rect 5813 47039 5871 47045
rect 5813 47005 5825 47039
rect 5859 47036 5871 47039
rect 6104 47036 6132 47076
rect 6178 47064 6184 47076
rect 6236 47104 6242 47116
rect 7285 47107 7343 47113
rect 7285 47104 7297 47107
rect 6236 47076 7297 47104
rect 6236 47064 6242 47076
rect 7285 47073 7297 47076
rect 7331 47073 7343 47107
rect 7285 47067 7343 47073
rect 7374 47064 7380 47116
rect 7432 47064 7438 47116
rect 5859 47008 6132 47036
rect 6273 47039 6331 47045
rect 5859 47005 5871 47008
rect 5813 46999 5871 47005
rect 6273 47005 6285 47039
rect 6319 47036 6331 47039
rect 6454 47036 6460 47048
rect 6319 47008 6460 47036
rect 6319 47005 6331 47008
rect 6273 46999 6331 47005
rect 6454 46996 6460 47008
rect 6512 47036 6518 47048
rect 7098 47036 7104 47048
rect 6512 47008 7104 47036
rect 6512 46996 6518 47008
rect 7098 46996 7104 47008
rect 7156 46996 7162 47048
rect 7193 47039 7251 47045
rect 7193 47005 7205 47039
rect 7239 47036 7251 47039
rect 8205 47039 8263 47045
rect 8205 47036 8217 47039
rect 7239 47008 8217 47036
rect 7239 47005 7251 47008
rect 7193 46999 7251 47005
rect 8205 47005 8217 47008
rect 8251 47036 8263 47039
rect 8864 47036 8892 47416
rect 8251 47008 8892 47036
rect 8251 47005 8263 47008
rect 8205 46999 8263 47005
rect 6086 46928 6092 46980
rect 6144 46968 6150 46980
rect 6641 46971 6699 46977
rect 6641 46968 6653 46971
rect 6144 46940 6653 46968
rect 6144 46928 6150 46940
rect 6641 46937 6653 46940
rect 6687 46937 6699 46971
rect 6641 46931 6699 46937
rect 5442 46860 5448 46912
rect 5500 46860 5506 46912
rect 5905 46903 5963 46909
rect 5905 46869 5917 46903
rect 5951 46900 5963 46903
rect 6178 46900 6184 46912
rect 5951 46872 6184 46900
rect 5951 46869 5963 46872
rect 5905 46863 5963 46869
rect 6178 46860 6184 46872
rect 6236 46860 6242 46912
rect 1104 46810 8832 46832
rect 1104 46758 3010 46810
rect 3062 46758 3074 46810
rect 3126 46758 3138 46810
rect 3190 46758 3202 46810
rect 3254 46758 3266 46810
rect 3318 46758 8010 46810
rect 8062 46758 8074 46810
rect 8126 46758 8138 46810
rect 8190 46758 8202 46810
rect 8254 46758 8266 46810
rect 8318 46758 8832 46810
rect 1104 46736 8832 46758
rect 6454 46628 6460 46640
rect 5934 46600 6460 46628
rect 6454 46588 6460 46600
rect 6512 46628 6518 46640
rect 8018 46628 8024 46640
rect 6512 46600 8024 46628
rect 6512 46588 6518 46600
rect 8018 46588 8024 46600
rect 8076 46588 8082 46640
rect 7193 46563 7251 46569
rect 7193 46529 7205 46563
rect 7239 46560 7251 46563
rect 8205 46563 8263 46569
rect 8205 46560 8217 46563
rect 7239 46532 8217 46560
rect 7239 46529 7251 46532
rect 7193 46523 7251 46529
rect 8205 46529 8217 46532
rect 8251 46560 8263 46563
rect 8251 46532 8616 46560
rect 8251 46529 8263 46532
rect 8205 46523 8263 46529
rect 4430 46452 4436 46504
rect 4488 46452 4494 46504
rect 4706 46452 4712 46504
rect 4764 46452 4770 46504
rect 6178 46452 6184 46504
rect 6236 46492 6242 46504
rect 7285 46495 7343 46501
rect 7285 46492 7297 46495
rect 6236 46464 7297 46492
rect 6236 46452 6242 46464
rect 7285 46461 7297 46464
rect 7331 46461 7343 46495
rect 7285 46455 7343 46461
rect 7374 46452 7380 46504
rect 7432 46492 7438 46504
rect 7834 46492 7840 46504
rect 7432 46464 7840 46492
rect 7432 46452 7438 46464
rect 7834 46452 7840 46464
rect 7892 46452 7898 46504
rect 6822 46316 6828 46368
rect 6880 46316 6886 46368
rect 8386 46316 8392 46368
rect 8444 46316 8450 46368
rect 8588 46356 8616 46532
rect 8588 46328 8892 46356
rect 1104 46266 8832 46288
rect 1104 46214 2350 46266
rect 2402 46214 2414 46266
rect 2466 46214 2478 46266
rect 2530 46214 2542 46266
rect 2594 46214 2606 46266
rect 2658 46214 7350 46266
rect 7402 46214 7414 46266
rect 7466 46214 7478 46266
rect 7530 46214 7542 46266
rect 7594 46214 7606 46266
rect 7658 46214 8832 46266
rect 1104 46192 8832 46214
rect 4706 46112 4712 46164
rect 4764 46152 4770 46164
rect 5169 46155 5227 46161
rect 5169 46152 5181 46155
rect 4764 46124 5181 46152
rect 4764 46112 4770 46124
rect 5169 46121 5181 46124
rect 5215 46121 5227 46155
rect 5169 46115 5227 46121
rect 6822 46112 6828 46164
rect 6880 46112 6886 46164
rect 8481 46155 8539 46161
rect 8481 46121 8493 46155
rect 8527 46152 8539 46155
rect 8864 46152 8892 46328
rect 8527 46124 8892 46152
rect 8527 46121 8539 46124
rect 8481 46115 8539 46121
rect 5994 45976 6000 46028
rect 6052 46016 6058 46028
rect 6089 46019 6147 46025
rect 6089 46016 6101 46019
rect 6052 45988 6101 46016
rect 6052 45976 6058 45988
rect 6089 45985 6101 45988
rect 6135 45985 6147 46019
rect 6840 46016 6868 46112
rect 6089 45979 6147 45985
rect 6472 45988 6868 46016
rect 5353 45951 5411 45957
rect 5353 45917 5365 45951
rect 5399 45948 5411 45951
rect 5442 45948 5448 45960
rect 5399 45920 5448 45948
rect 5399 45917 5411 45920
rect 5353 45911 5411 45917
rect 5442 45908 5448 45920
rect 5500 45908 5506 45960
rect 5905 45951 5963 45957
rect 5905 45917 5917 45951
rect 5951 45948 5963 45951
rect 6178 45948 6184 45960
rect 5951 45920 6184 45948
rect 5951 45917 5963 45920
rect 5905 45911 5963 45917
rect 6178 45908 6184 45920
rect 6236 45908 6242 45960
rect 6472 45957 6500 45988
rect 6457 45951 6515 45957
rect 6457 45917 6469 45951
rect 6503 45917 6515 45951
rect 6457 45911 6515 45917
rect 6546 45908 6552 45960
rect 6604 45948 6610 45960
rect 6733 45951 6791 45957
rect 6733 45948 6745 45951
rect 6604 45920 6745 45948
rect 6604 45908 6610 45920
rect 6733 45917 6745 45920
rect 6779 45917 6791 45951
rect 6733 45911 6791 45917
rect 8018 45908 8024 45960
rect 8076 45948 8082 45960
rect 8076 45920 8142 45948
rect 8076 45908 8082 45920
rect 7009 45883 7067 45889
rect 7009 45880 7021 45883
rect 6656 45852 7021 45880
rect 5537 45815 5595 45821
rect 5537 45781 5549 45815
rect 5583 45812 5595 45815
rect 5626 45812 5632 45824
rect 5583 45784 5632 45812
rect 5583 45781 5595 45784
rect 5537 45775 5595 45781
rect 5626 45772 5632 45784
rect 5684 45772 5690 45824
rect 5718 45772 5724 45824
rect 5776 45812 5782 45824
rect 5997 45815 6055 45821
rect 5997 45812 6009 45815
rect 5776 45784 6009 45812
rect 5776 45772 5782 45784
rect 5997 45781 6009 45784
rect 6043 45812 6055 45815
rect 6086 45812 6092 45824
rect 6043 45784 6092 45812
rect 6043 45781 6055 45784
rect 5997 45775 6055 45781
rect 6086 45772 6092 45784
rect 6144 45772 6150 45824
rect 6656 45821 6684 45852
rect 7009 45849 7021 45852
rect 7055 45849 7067 45883
rect 7009 45843 7067 45849
rect 6641 45815 6699 45821
rect 6641 45781 6653 45815
rect 6687 45781 6699 45815
rect 6641 45775 6699 45781
rect 1104 45722 8832 45744
rect 1104 45670 3010 45722
rect 3062 45670 3074 45722
rect 3126 45670 3138 45722
rect 3190 45670 3202 45722
rect 3254 45670 3266 45722
rect 3318 45670 8010 45722
rect 8062 45670 8074 45722
rect 8126 45670 8138 45722
rect 8190 45670 8202 45722
rect 8254 45670 8266 45722
rect 8318 45670 8832 45722
rect 1104 45648 8832 45670
rect 6086 45568 6092 45620
rect 6144 45568 6150 45620
rect 7285 45611 7343 45617
rect 7285 45577 7297 45611
rect 7331 45608 7343 45611
rect 7331 45580 7512 45608
rect 7331 45577 7343 45580
rect 7285 45571 7343 45577
rect 6104 45540 6132 45568
rect 7377 45543 7435 45549
rect 7377 45540 7389 45543
rect 6104 45512 7389 45540
rect 7377 45509 7389 45512
rect 7423 45509 7435 45543
rect 7484 45540 7512 45580
rect 7484 45512 8800 45540
rect 7377 45503 7435 45509
rect 6454 45472 6460 45484
rect 5750 45444 6460 45472
rect 6454 45432 6460 45444
rect 6512 45432 6518 45484
rect 6914 45432 6920 45484
rect 6972 45472 6978 45484
rect 7098 45472 7104 45484
rect 6972 45444 7104 45472
rect 6972 45432 6978 45444
rect 7098 45432 7104 45444
rect 7156 45472 7162 45484
rect 7745 45475 7803 45481
rect 7745 45472 7757 45475
rect 7156 45444 7757 45472
rect 7156 45432 7162 45444
rect 7745 45441 7757 45444
rect 7791 45441 7803 45475
rect 7745 45435 7803 45441
rect 4341 45407 4399 45413
rect 4341 45373 4353 45407
rect 4387 45404 4399 45407
rect 4387 45376 4476 45404
rect 4387 45373 4399 45376
rect 4341 45367 4399 45373
rect 4448 45280 4476 45376
rect 4614 45364 4620 45416
rect 4672 45364 4678 45416
rect 7561 45407 7619 45413
rect 7561 45373 7573 45407
rect 7607 45404 7619 45407
rect 7834 45404 7840 45416
rect 7607 45376 7840 45404
rect 7607 45373 7619 45376
rect 7561 45367 7619 45373
rect 7834 45364 7840 45376
rect 7892 45404 7898 45416
rect 7929 45407 7987 45413
rect 7929 45404 7941 45407
rect 7892 45376 7941 45404
rect 7892 45364 7898 45376
rect 7929 45373 7941 45376
rect 7975 45373 7987 45407
rect 7929 45367 7987 45373
rect 4430 45228 4436 45280
rect 4488 45228 4494 45280
rect 6914 45228 6920 45280
rect 6972 45228 6978 45280
rect 8772 45268 8800 45512
rect 8772 45240 8892 45268
rect 1104 45178 8832 45200
rect 1104 45126 2350 45178
rect 2402 45126 2414 45178
rect 2466 45126 2478 45178
rect 2530 45126 2542 45178
rect 2594 45126 2606 45178
rect 2658 45126 7350 45178
rect 7402 45126 7414 45178
rect 7466 45126 7478 45178
rect 7530 45126 7542 45178
rect 7594 45126 7606 45178
rect 7658 45126 8832 45178
rect 1104 45104 8832 45126
rect 4614 45024 4620 45076
rect 4672 45064 4678 45076
rect 5261 45067 5319 45073
rect 5261 45064 5273 45067
rect 4672 45036 5273 45064
rect 4672 45024 4678 45036
rect 5261 45033 5273 45036
rect 5307 45033 5319 45067
rect 5261 45027 5319 45033
rect 8481 45067 8539 45073
rect 8481 45033 8493 45067
rect 8527 45064 8539 45067
rect 8864 45064 8892 45240
rect 8527 45036 8892 45064
rect 8527 45033 8539 45036
rect 8481 45027 8539 45033
rect 5445 44863 5503 44869
rect 5445 44829 5457 44863
rect 5491 44860 5503 44863
rect 5626 44860 5632 44872
rect 5491 44832 5632 44860
rect 5491 44829 5503 44832
rect 5445 44823 5503 44829
rect 5626 44820 5632 44832
rect 5684 44820 5690 44872
rect 6546 44820 6552 44872
rect 6604 44860 6610 44872
rect 6733 44863 6791 44869
rect 6733 44860 6745 44863
rect 6604 44832 6745 44860
rect 6604 44820 6610 44832
rect 6733 44829 6745 44832
rect 6779 44829 6791 44863
rect 6733 44823 6791 44829
rect 8018 44820 8024 44872
rect 8076 44860 8082 44872
rect 8076 44832 8142 44860
rect 8076 44820 8082 44832
rect 7009 44795 7067 44801
rect 7009 44761 7021 44795
rect 7055 44761 7067 44795
rect 7009 44755 7067 44761
rect 7024 44724 7052 44755
rect 7190 44724 7196 44736
rect 7024 44696 7196 44724
rect 7190 44684 7196 44696
rect 7248 44684 7254 44736
rect 1104 44634 8832 44656
rect 1104 44582 3010 44634
rect 3062 44582 3074 44634
rect 3126 44582 3138 44634
rect 3190 44582 3202 44634
rect 3254 44582 3266 44634
rect 3318 44582 8010 44634
rect 8062 44582 8074 44634
rect 8126 44582 8138 44634
rect 8190 44582 8202 44634
rect 8254 44582 8266 44634
rect 8318 44582 8832 44634
rect 1104 44560 8832 44582
rect 6914 44480 6920 44532
rect 6972 44480 6978 44532
rect 7009 44523 7067 44529
rect 7009 44489 7021 44523
rect 7055 44520 7067 44523
rect 7190 44520 7196 44532
rect 7055 44492 7196 44520
rect 7055 44489 7067 44492
rect 7009 44483 7067 44489
rect 7190 44480 7196 44492
rect 7248 44480 7254 44532
rect 8386 44480 8392 44532
rect 8444 44480 8450 44532
rect 5350 44344 5356 44396
rect 5408 44344 5414 44396
rect 6932 44384 6960 44480
rect 7193 44387 7251 44393
rect 7193 44384 7205 44387
rect 6932 44356 7205 44384
rect 7193 44353 7205 44356
rect 7239 44353 7251 44387
rect 7193 44347 7251 44353
rect 8205 44387 8263 44393
rect 8205 44353 8217 44387
rect 8251 44384 8263 44387
rect 8864 44384 8892 45036
rect 8251 44356 8892 44384
rect 8251 44353 8263 44356
rect 8205 44347 8263 44353
rect 5166 44140 5172 44192
rect 5224 44140 5230 44192
rect 1104 44090 8832 44112
rect 1104 44038 2350 44090
rect 2402 44038 2414 44090
rect 2466 44038 2478 44090
rect 2530 44038 2542 44090
rect 2594 44038 2606 44090
rect 2658 44038 7350 44090
rect 7402 44038 7414 44090
rect 7466 44038 7478 44090
rect 7530 44038 7542 44090
rect 7594 44038 7606 44090
rect 7658 44038 8832 44090
rect 1104 44016 8832 44038
rect 6270 43936 6276 43988
rect 6328 43976 6334 43988
rect 6641 43979 6699 43985
rect 6641 43976 6653 43979
rect 6328 43948 6653 43976
rect 6328 43936 6334 43948
rect 6641 43945 6653 43948
rect 6687 43945 6699 43979
rect 6641 43939 6699 43945
rect 5166 43800 5172 43852
rect 5224 43800 5230 43852
rect 4430 43732 4436 43784
rect 4488 43772 4494 43784
rect 4893 43775 4951 43781
rect 4893 43772 4905 43775
rect 4488 43744 4905 43772
rect 4488 43732 4494 43744
rect 4893 43741 4905 43744
rect 4939 43741 4951 43775
rect 6454 43772 6460 43784
rect 6302 43744 6460 43772
rect 4893 43735 4951 43741
rect 6454 43732 6460 43744
rect 6512 43732 6518 43784
rect 8481 43775 8539 43781
rect 8481 43741 8493 43775
rect 8527 43772 8539 43775
rect 8527 43744 8892 43772
rect 8527 43741 8539 43744
rect 8481 43735 8539 43741
rect 8864 43648 8892 43744
rect 7926 43596 7932 43648
rect 7984 43636 7990 43648
rect 8297 43639 8355 43645
rect 8297 43636 8309 43639
rect 7984 43608 8309 43636
rect 7984 43596 7990 43608
rect 8297 43605 8309 43608
rect 8343 43605 8355 43639
rect 8297 43599 8355 43605
rect 8846 43596 8852 43648
rect 8904 43596 8910 43648
rect 1104 43546 8832 43568
rect 1104 43494 3010 43546
rect 3062 43494 3074 43546
rect 3126 43494 3138 43546
rect 3190 43494 3202 43546
rect 3254 43494 3266 43546
rect 3318 43494 8010 43546
rect 8062 43494 8074 43546
rect 8126 43494 8138 43546
rect 8190 43494 8202 43546
rect 8254 43494 8266 43546
rect 8318 43494 8832 43546
rect 1104 43472 8832 43494
rect 5350 43392 5356 43444
rect 5408 43392 5414 43444
rect 5813 43435 5871 43441
rect 5813 43401 5825 43435
rect 5859 43432 5871 43435
rect 6270 43432 6276 43444
rect 5859 43404 6276 43432
rect 5859 43401 5871 43404
rect 5813 43395 5871 43401
rect 6270 43392 6276 43404
rect 6328 43392 6334 43444
rect 6733 43435 6791 43441
rect 6733 43401 6745 43435
rect 6779 43432 6791 43435
rect 6914 43432 6920 43444
rect 6779 43404 6920 43432
rect 6779 43401 6791 43404
rect 6733 43395 6791 43401
rect 6914 43392 6920 43404
rect 6972 43432 6978 43444
rect 7098 43432 7104 43444
rect 6972 43404 7104 43432
rect 6972 43392 6978 43404
rect 7098 43392 7104 43404
rect 7156 43392 7162 43444
rect 5721 43299 5779 43305
rect 5721 43265 5733 43299
rect 5767 43296 5779 43299
rect 6178 43296 6184 43308
rect 5767 43268 6184 43296
rect 5767 43265 5779 43268
rect 5721 43259 5779 43265
rect 6178 43256 6184 43268
rect 6236 43256 6242 43308
rect 6917 43299 6975 43305
rect 6917 43265 6929 43299
rect 6963 43296 6975 43299
rect 7098 43296 7104 43308
rect 6963 43268 7104 43296
rect 6963 43265 6975 43268
rect 6917 43259 6975 43265
rect 7098 43256 7104 43268
rect 7156 43256 7162 43308
rect 7190 43256 7196 43308
rect 7248 43296 7254 43308
rect 7285 43299 7343 43305
rect 7285 43296 7297 43299
rect 7248 43268 7297 43296
rect 7248 43256 7254 43268
rect 7285 43265 7297 43268
rect 7331 43265 7343 43299
rect 7285 43259 7343 43265
rect 5994 43188 6000 43240
rect 6052 43228 6058 43240
rect 6457 43231 6515 43237
rect 6457 43228 6469 43231
rect 6052 43200 6469 43228
rect 6052 43188 6058 43200
rect 6457 43197 6469 43200
rect 6503 43197 6515 43231
rect 6457 43191 6515 43197
rect 6914 43052 6920 43104
rect 6972 43092 6978 43104
rect 7101 43095 7159 43101
rect 7101 43092 7113 43095
rect 6972 43064 7113 43092
rect 6972 43052 6978 43064
rect 7101 43061 7113 43064
rect 7147 43061 7159 43095
rect 7101 43055 7159 43061
rect 1104 43002 8832 43024
rect 1104 42950 2350 43002
rect 2402 42950 2414 43002
rect 2466 42950 2478 43002
rect 2530 42950 2542 43002
rect 2594 42950 2606 43002
rect 2658 42950 7350 43002
rect 7402 42950 7414 43002
rect 7466 42950 7478 43002
rect 7530 42950 7542 43002
rect 7594 42950 7606 43002
rect 7658 42950 8832 43002
rect 1104 42928 8832 42950
rect 6812 42891 6870 42897
rect 6812 42857 6824 42891
rect 6858 42888 6870 42891
rect 6914 42888 6920 42900
rect 6858 42860 6920 42888
rect 6858 42857 6870 42860
rect 6812 42851 6870 42857
rect 6914 42848 6920 42860
rect 6972 42848 6978 42900
rect 6546 42712 6552 42764
rect 6604 42712 6610 42764
rect 4430 42644 4436 42696
rect 4488 42684 4494 42696
rect 4709 42687 4767 42693
rect 4709 42684 4721 42687
rect 4488 42656 4721 42684
rect 4488 42644 4494 42656
rect 4709 42653 4721 42656
rect 4755 42653 4767 42687
rect 6454 42684 6460 42696
rect 6118 42656 6460 42684
rect 4709 42647 4767 42653
rect 6454 42644 6460 42656
rect 6512 42644 6518 42696
rect 4982 42576 4988 42628
rect 5040 42576 5046 42628
rect 6472 42616 6500 42644
rect 6822 42616 6828 42628
rect 6472 42588 6828 42616
rect 6822 42576 6828 42588
rect 6880 42616 6886 42628
rect 6880 42588 7314 42616
rect 6880 42576 6886 42588
rect 6457 42551 6515 42557
rect 6457 42517 6469 42551
rect 6503 42548 6515 42551
rect 7098 42548 7104 42560
rect 6503 42520 7104 42548
rect 6503 42517 6515 42520
rect 6457 42511 6515 42517
rect 7098 42508 7104 42520
rect 7156 42508 7162 42560
rect 7834 42508 7840 42560
rect 7892 42548 7898 42560
rect 8297 42551 8355 42557
rect 8297 42548 8309 42551
rect 7892 42520 8309 42548
rect 7892 42508 7898 42520
rect 8297 42517 8309 42520
rect 8343 42517 8355 42551
rect 8297 42511 8355 42517
rect 1104 42458 8832 42480
rect 1104 42406 3010 42458
rect 3062 42406 3074 42458
rect 3126 42406 3138 42458
rect 3190 42406 3202 42458
rect 3254 42406 3266 42458
rect 3318 42406 8010 42458
rect 8062 42406 8074 42458
rect 8126 42406 8138 42458
rect 8190 42406 8202 42458
rect 8254 42406 8266 42458
rect 8318 42406 8832 42458
rect 1104 42384 8832 42406
rect 4982 42304 4988 42356
rect 5040 42344 5046 42356
rect 5261 42347 5319 42353
rect 5261 42344 5273 42347
rect 5040 42316 5273 42344
rect 5040 42304 5046 42316
rect 5261 42313 5273 42316
rect 5307 42313 5319 42347
rect 7098 42344 7104 42356
rect 5261 42307 5319 42313
rect 6012 42316 7104 42344
rect 5813 42279 5871 42285
rect 5813 42245 5825 42279
rect 5859 42276 5871 42279
rect 5902 42276 5908 42288
rect 5859 42248 5908 42276
rect 5859 42245 5871 42248
rect 5813 42239 5871 42245
rect 5902 42236 5908 42248
rect 5960 42236 5966 42288
rect 6012 42285 6040 42316
rect 7098 42304 7104 42316
rect 7156 42304 7162 42356
rect 7190 42304 7196 42356
rect 7248 42344 7254 42356
rect 7285 42347 7343 42353
rect 7285 42344 7297 42347
rect 7248 42316 7297 42344
rect 7248 42304 7254 42316
rect 7285 42313 7297 42316
rect 7331 42313 7343 42347
rect 7285 42307 7343 42313
rect 7653 42347 7711 42353
rect 7653 42313 7665 42347
rect 7699 42344 7711 42347
rect 8021 42347 8079 42353
rect 8021 42344 8033 42347
rect 7699 42316 8033 42344
rect 7699 42313 7711 42316
rect 7653 42307 7711 42313
rect 8021 42313 8033 42316
rect 8067 42313 8079 42347
rect 8021 42307 8079 42313
rect 5997 42279 6055 42285
rect 5997 42245 6009 42279
rect 6043 42245 6055 42279
rect 5997 42239 6055 42245
rect 6178 42236 6184 42288
rect 6236 42276 6242 42288
rect 6825 42279 6883 42285
rect 6825 42276 6837 42279
rect 6236 42248 6837 42276
rect 6236 42236 6242 42248
rect 6825 42245 6837 42248
rect 6871 42245 6883 42279
rect 6825 42239 6883 42245
rect 6917 42279 6975 42285
rect 6917 42245 6929 42279
rect 6963 42276 6975 42279
rect 7834 42276 7840 42288
rect 6963 42248 7840 42276
rect 6963 42245 6975 42248
rect 6917 42239 6975 42245
rect 7834 42236 7840 42248
rect 7892 42236 7898 42288
rect 7926 42236 7932 42288
rect 7984 42276 7990 42288
rect 8113 42279 8171 42285
rect 8113 42276 8125 42279
rect 7984 42248 8125 42276
rect 7984 42236 7990 42248
rect 8113 42245 8125 42248
rect 8159 42245 8171 42279
rect 8113 42239 8171 42245
rect 5445 42211 5503 42217
rect 5445 42177 5457 42211
rect 5491 42208 5503 42211
rect 5629 42211 5687 42217
rect 5629 42208 5641 42211
rect 5491 42180 5641 42208
rect 5491 42177 5503 42180
rect 5445 42171 5503 42177
rect 5629 42177 5641 42180
rect 5675 42177 5687 42211
rect 5629 42171 5687 42177
rect 7469 42211 7527 42217
rect 7469 42177 7481 42211
rect 7515 42177 7527 42211
rect 7469 42171 7527 42177
rect 6733 42143 6791 42149
rect 6733 42109 6745 42143
rect 6779 42140 6791 42143
rect 6914 42140 6920 42152
rect 6779 42112 6920 42140
rect 6779 42109 6791 42112
rect 6733 42103 6791 42109
rect 6914 42100 6920 42112
rect 6972 42100 6978 42152
rect 7484 42072 7512 42171
rect 7852 42149 7880 42236
rect 7837 42143 7895 42149
rect 7837 42109 7849 42143
rect 7883 42109 7895 42143
rect 7837 42103 7895 42109
rect 8386 42072 8392 42084
rect 7484 42044 8392 42072
rect 8386 42032 8392 42044
rect 8444 42032 8450 42084
rect 8481 42007 8539 42013
rect 8481 41973 8493 42007
rect 8527 42004 8539 42007
rect 8527 41976 8892 42004
rect 8527 41973 8539 41976
rect 8481 41967 8539 41973
rect 1104 41914 8832 41936
rect 1104 41862 2350 41914
rect 2402 41862 2414 41914
rect 2466 41862 2478 41914
rect 2530 41862 2542 41914
rect 2594 41862 2606 41914
rect 2658 41862 7350 41914
rect 7402 41862 7414 41914
rect 7466 41862 7478 41914
rect 7530 41862 7542 41914
rect 7594 41862 7606 41914
rect 7658 41862 8832 41914
rect 1104 41840 8832 41862
rect 5902 41760 5908 41812
rect 5960 41800 5966 41812
rect 6549 41803 6607 41809
rect 6549 41800 6561 41803
rect 5960 41772 6561 41800
rect 5960 41760 5966 41772
rect 6549 41769 6561 41772
rect 6595 41769 6607 41803
rect 6549 41763 6607 41769
rect 5813 41599 5871 41605
rect 5813 41565 5825 41599
rect 5859 41596 5871 41599
rect 6457 41599 6515 41605
rect 6457 41596 6469 41599
rect 5859 41568 6469 41596
rect 5859 41565 5871 41568
rect 5813 41559 5871 41565
rect 6457 41565 6469 41568
rect 6503 41596 6515 41599
rect 6730 41596 6736 41608
rect 6503 41568 6736 41596
rect 6503 41565 6515 41568
rect 6457 41559 6515 41565
rect 6730 41556 6736 41568
rect 6788 41556 6794 41608
rect 6914 41556 6920 41608
rect 6972 41596 6978 41608
rect 7469 41599 7527 41605
rect 7469 41596 7481 41599
rect 6972 41568 7481 41596
rect 6972 41556 6978 41568
rect 7469 41565 7481 41568
rect 7515 41565 7527 41599
rect 7469 41559 7527 41565
rect 8205 41599 8263 41605
rect 8205 41565 8217 41599
rect 8251 41596 8263 41599
rect 8864 41596 8892 41976
rect 8251 41568 8892 41596
rect 8251 41565 8263 41568
rect 8205 41559 8263 41565
rect 6178 41488 6184 41540
rect 6236 41488 6242 41540
rect 7834 41488 7840 41540
rect 7892 41528 7898 41540
rect 8021 41531 8079 41537
rect 8021 41528 8033 41531
rect 7892 41500 8033 41528
rect 7892 41488 7898 41500
rect 8021 41497 8033 41500
rect 8067 41497 8079 41531
rect 8021 41491 8079 41497
rect 7377 41463 7435 41469
rect 7377 41429 7389 41463
rect 7423 41460 7435 41463
rect 7742 41460 7748 41472
rect 7423 41432 7748 41460
rect 7423 41429 7435 41432
rect 7377 41423 7435 41429
rect 7742 41420 7748 41432
rect 7800 41420 7806 41472
rect 1104 41370 8832 41392
rect 1104 41318 3010 41370
rect 3062 41318 3074 41370
rect 3126 41318 3138 41370
rect 3190 41318 3202 41370
rect 3254 41318 3266 41370
rect 3318 41318 8010 41370
rect 8062 41318 8074 41370
rect 8126 41318 8138 41370
rect 8190 41318 8202 41370
rect 8254 41318 8266 41370
rect 8318 41318 8832 41370
rect 1104 41296 8832 41318
rect 6086 41216 6092 41268
rect 6144 41256 6150 41268
rect 6181 41259 6239 41265
rect 6181 41256 6193 41259
rect 6144 41228 6193 41256
rect 6144 41216 6150 41228
rect 6181 41225 6193 41228
rect 6227 41225 6239 41259
rect 6181 41219 6239 41225
rect 6914 41188 6920 41200
rect 5934 41160 6920 41188
rect 6914 41148 6920 41160
rect 6972 41188 6978 41200
rect 7098 41188 7104 41200
rect 6972 41160 7104 41188
rect 6972 41148 6978 41160
rect 7098 41148 7104 41160
rect 7156 41148 7162 41200
rect 4430 41080 4436 41132
rect 4488 41080 4494 41132
rect 6454 41080 6460 41132
rect 6512 41080 6518 41132
rect 8205 41123 8263 41129
rect 8205 41089 8217 41123
rect 8251 41120 8263 41123
rect 8251 41092 8892 41120
rect 8251 41089 8263 41092
rect 8205 41083 8263 41089
rect 4706 41012 4712 41064
rect 4764 41012 4770 41064
rect 6641 40919 6699 40925
rect 6641 40885 6653 40919
rect 6687 40916 6699 40919
rect 6914 40916 6920 40928
rect 6687 40888 6920 40916
rect 6687 40885 6699 40888
rect 6641 40879 6699 40885
rect 6914 40876 6920 40888
rect 6972 40876 6978 40928
rect 8386 40876 8392 40928
rect 8444 40876 8450 40928
rect 1104 40826 8832 40848
rect 1104 40774 2350 40826
rect 2402 40774 2414 40826
rect 2466 40774 2478 40826
rect 2530 40774 2542 40826
rect 2594 40774 2606 40826
rect 2658 40774 7350 40826
rect 7402 40774 7414 40826
rect 7466 40774 7478 40826
rect 7530 40774 7542 40826
rect 7594 40774 7606 40826
rect 7658 40774 8832 40826
rect 1104 40752 8832 40774
rect 4617 40715 4675 40721
rect 4617 40681 4629 40715
rect 4663 40712 4675 40715
rect 4706 40712 4712 40724
rect 4663 40684 4712 40712
rect 4663 40681 4675 40684
rect 4617 40675 4675 40681
rect 4706 40672 4712 40684
rect 4764 40672 4770 40724
rect 7006 40576 7012 40588
rect 6656 40548 7012 40576
rect 4798 40468 4804 40520
rect 4856 40468 4862 40520
rect 6656 40517 6684 40548
rect 7006 40536 7012 40548
rect 7064 40536 7070 40588
rect 6641 40511 6699 40517
rect 6641 40477 6653 40511
rect 6687 40477 6699 40511
rect 6641 40471 6699 40477
rect 6730 40468 6736 40520
rect 6788 40468 6794 40520
rect 6914 40400 6920 40452
rect 6972 40440 6978 40452
rect 7009 40443 7067 40449
rect 7009 40440 7021 40443
rect 6972 40412 7021 40440
rect 6972 40400 6978 40412
rect 7009 40409 7021 40412
rect 7055 40409 7067 40443
rect 7009 40403 7067 40409
rect 7098 40400 7104 40452
rect 7156 40440 7162 40452
rect 7156 40412 7498 40440
rect 7156 40400 7162 40412
rect 5353 40375 5411 40381
rect 5353 40341 5365 40375
rect 5399 40372 5411 40375
rect 5534 40372 5540 40384
rect 5399 40344 5540 40372
rect 5399 40341 5411 40344
rect 5353 40335 5411 40341
rect 5534 40332 5540 40344
rect 5592 40372 5598 40384
rect 6822 40372 6828 40384
rect 5592 40344 6828 40372
rect 5592 40332 5598 40344
rect 6822 40332 6828 40344
rect 6880 40332 6886 40384
rect 8481 40375 8539 40381
rect 8481 40341 8493 40375
rect 8527 40372 8539 40375
rect 8864 40372 8892 41092
rect 8527 40344 8892 40372
rect 8527 40341 8539 40344
rect 8481 40335 8539 40341
rect 1104 40282 8832 40304
rect 1104 40230 3010 40282
rect 3062 40230 3074 40282
rect 3126 40230 3138 40282
rect 3190 40230 3202 40282
rect 3254 40230 3266 40282
rect 3318 40230 8010 40282
rect 8062 40230 8074 40282
rect 8126 40230 8138 40282
rect 8190 40230 8202 40282
rect 8254 40230 8266 40282
rect 8318 40230 8832 40282
rect 1104 40208 8832 40230
rect 4798 40128 4804 40180
rect 4856 40168 4862 40180
rect 5261 40171 5319 40177
rect 5261 40168 5273 40171
rect 4856 40140 5273 40168
rect 4856 40128 4862 40140
rect 5261 40137 5273 40140
rect 5307 40137 5319 40171
rect 5261 40131 5319 40137
rect 5721 40171 5779 40177
rect 5721 40137 5733 40171
rect 5767 40168 5779 40171
rect 6086 40168 6092 40180
rect 5767 40140 6092 40168
rect 5767 40137 5779 40140
rect 5721 40131 5779 40137
rect 6086 40128 6092 40140
rect 6144 40128 6150 40180
rect 6362 40128 6368 40180
rect 6420 40128 6426 40180
rect 6454 40128 6460 40180
rect 6512 40168 6518 40180
rect 6733 40171 6791 40177
rect 6733 40168 6745 40171
rect 6512 40140 6745 40168
rect 6512 40128 6518 40140
rect 6733 40137 6745 40140
rect 6779 40137 6791 40171
rect 6733 40131 6791 40137
rect 7101 40171 7159 40177
rect 7101 40137 7113 40171
rect 7147 40168 7159 40171
rect 8864 40168 8892 40344
rect 7147 40140 8892 40168
rect 7147 40137 7159 40140
rect 7101 40131 7159 40137
rect 5626 40060 5632 40112
rect 5684 40060 5690 40112
rect 6380 40041 6408 40128
rect 6365 40035 6423 40041
rect 6365 40001 6377 40035
rect 6411 40001 6423 40035
rect 6365 39995 6423 40001
rect 5902 39924 5908 39976
rect 5960 39924 5966 39976
rect 6270 39924 6276 39976
rect 6328 39964 6334 39976
rect 7193 39967 7251 39973
rect 7193 39964 7205 39967
rect 6328 39936 7205 39964
rect 6328 39924 6334 39936
rect 7193 39933 7205 39936
rect 7239 39933 7251 39967
rect 7193 39927 7251 39933
rect 7377 39967 7435 39973
rect 7377 39933 7389 39967
rect 7423 39964 7435 39967
rect 7742 39964 7748 39976
rect 7423 39936 7748 39964
rect 7423 39933 7435 39936
rect 7377 39927 7435 39933
rect 7742 39924 7748 39936
rect 7800 39924 7806 39976
rect 6546 39788 6552 39840
rect 6604 39788 6610 39840
rect 1104 39738 8832 39760
rect 1104 39686 2350 39738
rect 2402 39686 2414 39738
rect 2466 39686 2478 39738
rect 2530 39686 2542 39738
rect 2594 39686 2606 39738
rect 2658 39686 7350 39738
rect 7402 39686 7414 39738
rect 7466 39686 7478 39738
rect 7530 39686 7542 39738
rect 7594 39686 7606 39738
rect 7658 39686 8832 39738
rect 1104 39664 8832 39686
rect 4430 39380 4436 39432
rect 4488 39420 4494 39432
rect 4709 39423 4767 39429
rect 4709 39420 4721 39423
rect 4488 39392 4721 39420
rect 4488 39380 4494 39392
rect 4709 39389 4721 39392
rect 4755 39389 4767 39423
rect 4709 39383 4767 39389
rect 6730 39380 6736 39432
rect 6788 39380 6794 39432
rect 4982 39312 4988 39364
rect 5040 39312 5046 39364
rect 6546 39352 6552 39364
rect 6210 39324 6552 39352
rect 6546 39312 6552 39324
rect 6604 39312 6610 39364
rect 7009 39355 7067 39361
rect 7009 39321 7021 39355
rect 7055 39321 7067 39355
rect 7009 39315 7067 39321
rect 5902 39244 5908 39296
rect 5960 39284 5966 39296
rect 6457 39287 6515 39293
rect 6457 39284 6469 39287
rect 5960 39256 6469 39284
rect 5960 39244 5966 39256
rect 6457 39253 6469 39256
rect 6503 39253 6515 39287
rect 7024 39284 7052 39315
rect 7098 39312 7104 39364
rect 7156 39352 7162 39364
rect 7156 39324 7498 39352
rect 7156 39312 7162 39324
rect 7650 39284 7656 39296
rect 7024 39256 7656 39284
rect 6457 39247 6515 39253
rect 7650 39244 7656 39256
rect 7708 39244 7714 39296
rect 8481 39287 8539 39293
rect 8481 39253 8493 39287
rect 8527 39284 8539 39287
rect 8527 39256 8892 39284
rect 8527 39253 8539 39256
rect 8481 39247 8539 39253
rect 1104 39194 8832 39216
rect 1104 39142 3010 39194
rect 3062 39142 3074 39194
rect 3126 39142 3138 39194
rect 3190 39142 3202 39194
rect 3254 39142 3266 39194
rect 3318 39142 8010 39194
rect 8062 39142 8074 39194
rect 8126 39142 8138 39194
rect 8190 39142 8202 39194
rect 8254 39142 8266 39194
rect 8318 39142 8832 39194
rect 1104 39120 8832 39142
rect 4982 39040 4988 39092
rect 5040 39080 5046 39092
rect 5169 39083 5227 39089
rect 5169 39080 5181 39083
rect 5040 39052 5181 39080
rect 5040 39040 5046 39052
rect 5169 39049 5181 39052
rect 5215 39049 5227 39083
rect 5169 39043 5227 39049
rect 5445 39083 5503 39089
rect 5445 39049 5457 39083
rect 5491 39049 5503 39083
rect 5445 39043 5503 39049
rect 7469 39083 7527 39089
rect 7469 39049 7481 39083
rect 7515 39049 7527 39083
rect 7469 39043 7527 39049
rect 7561 39083 7619 39089
rect 7561 39049 7573 39083
rect 7607 39080 7619 39083
rect 7650 39080 7656 39092
rect 7607 39052 7656 39080
rect 7607 39049 7619 39052
rect 7561 39043 7619 39049
rect 5353 38947 5411 38953
rect 5353 38913 5365 38947
rect 5399 38944 5411 38947
rect 5460 38944 5488 39043
rect 5813 39015 5871 39021
rect 5813 38981 5825 39015
rect 5859 39012 5871 39015
rect 6270 39012 6276 39024
rect 5859 38984 6276 39012
rect 5859 38981 5871 38984
rect 5813 38975 5871 38981
rect 6270 38972 6276 38984
rect 6328 38972 6334 39024
rect 5399 38916 5488 38944
rect 5399 38913 5411 38916
rect 5353 38907 5411 38913
rect 5902 38904 5908 38956
rect 5960 38944 5966 38956
rect 7009 38947 7067 38953
rect 7009 38944 7021 38947
rect 5960 38916 7021 38944
rect 5960 38904 5966 38916
rect 7009 38913 7021 38916
rect 7055 38913 7067 38947
rect 7009 38907 7067 38913
rect 7101 38947 7159 38953
rect 7101 38913 7113 38947
rect 7147 38913 7159 38947
rect 7484 38944 7512 39043
rect 7650 39040 7656 39052
rect 7708 39040 7714 39092
rect 8386 39040 8392 39092
rect 8444 39040 8450 39092
rect 7745 38947 7803 38953
rect 7745 38944 7757 38947
rect 7484 38916 7757 38944
rect 7101 38907 7159 38913
rect 7745 38913 7757 38916
rect 7791 38913 7803 38947
rect 7745 38907 7803 38913
rect 8205 38947 8263 38953
rect 8205 38913 8217 38947
rect 8251 38944 8263 38947
rect 8864 38944 8892 39256
rect 8251 38916 8892 38944
rect 8251 38913 8263 38916
rect 8205 38907 8263 38913
rect 6086 38836 6092 38888
rect 6144 38836 6150 38888
rect 6917 38879 6975 38885
rect 6917 38845 6929 38879
rect 6963 38845 6975 38879
rect 7116 38876 7144 38907
rect 8220 38876 8248 38907
rect 7116 38848 8248 38876
rect 6917 38839 6975 38845
rect 6932 38808 6960 38839
rect 7190 38808 7196 38820
rect 6932 38780 7196 38808
rect 7190 38768 7196 38780
rect 7248 38808 7254 38820
rect 7742 38808 7748 38820
rect 7248 38780 7748 38808
rect 7248 38768 7254 38780
rect 7742 38768 7748 38780
rect 7800 38768 7806 38820
rect 1104 38650 8832 38672
rect 1104 38598 2350 38650
rect 2402 38598 2414 38650
rect 2466 38598 2478 38650
rect 2530 38598 2542 38650
rect 2594 38598 2606 38650
rect 2658 38598 7350 38650
rect 7402 38598 7414 38650
rect 7466 38598 7478 38650
rect 7530 38598 7542 38650
rect 7594 38598 7606 38650
rect 7658 38598 8832 38650
rect 1104 38576 8832 38598
rect 6733 38471 6791 38477
rect 6733 38437 6745 38471
rect 6779 38468 6791 38471
rect 6779 38440 6813 38468
rect 6779 38437 6791 38440
rect 6733 38431 6791 38437
rect 6748 38400 6776 38431
rect 7098 38400 7104 38412
rect 6012 38372 7104 38400
rect 6012 38344 6040 38372
rect 7098 38360 7104 38372
rect 7156 38360 7162 38412
rect 4430 38292 4436 38344
rect 4488 38332 4494 38344
rect 4617 38335 4675 38341
rect 4617 38332 4629 38335
rect 4488 38304 4629 38332
rect 4488 38292 4494 38304
rect 4617 38301 4629 38304
rect 4663 38301 4675 38335
rect 4617 38295 4675 38301
rect 5994 38292 6000 38344
rect 6052 38292 6058 38344
rect 7742 38292 7748 38344
rect 7800 38332 7806 38344
rect 8205 38335 8263 38341
rect 8205 38332 8217 38335
rect 7800 38304 8217 38332
rect 7800 38292 7806 38304
rect 8205 38301 8217 38304
rect 8251 38301 8263 38335
rect 8205 38295 8263 38301
rect 4890 38224 4896 38276
rect 4948 38224 4954 38276
rect 6546 38224 6552 38276
rect 6604 38224 6610 38276
rect 5810 38156 5816 38208
rect 5868 38196 5874 38208
rect 6365 38199 6423 38205
rect 6365 38196 6377 38199
rect 5868 38168 6377 38196
rect 5868 38156 5874 38168
rect 6365 38165 6377 38168
rect 6411 38165 6423 38199
rect 6365 38159 6423 38165
rect 8386 38156 8392 38208
rect 8444 38156 8450 38208
rect 1104 38106 8832 38128
rect 1104 38054 3010 38106
rect 3062 38054 3074 38106
rect 3126 38054 3138 38106
rect 3190 38054 3202 38106
rect 3254 38054 3266 38106
rect 3318 38054 8010 38106
rect 8062 38054 8074 38106
rect 8126 38054 8138 38106
rect 8190 38054 8202 38106
rect 8254 38054 8266 38106
rect 8318 38054 8832 38106
rect 1104 38032 8832 38054
rect 4890 37952 4896 38004
rect 4948 37992 4954 38004
rect 5077 37995 5135 38001
rect 5077 37992 5089 37995
rect 4948 37964 5089 37992
rect 4948 37952 4954 37964
rect 5077 37961 5089 37964
rect 5123 37961 5135 37995
rect 5077 37955 5135 37961
rect 5445 37995 5503 38001
rect 5445 37961 5457 37995
rect 5491 37961 5503 37995
rect 5445 37955 5503 37961
rect 5813 37995 5871 38001
rect 5813 37961 5825 37995
rect 5859 37992 5871 37995
rect 5902 37992 5908 38004
rect 5859 37964 5908 37992
rect 5859 37961 5871 37964
rect 5813 37955 5871 37961
rect 5261 37859 5319 37865
rect 5261 37825 5273 37859
rect 5307 37856 5319 37859
rect 5460 37856 5488 37955
rect 5902 37952 5908 37964
rect 5960 37952 5966 38004
rect 6641 37995 6699 38001
rect 6641 37961 6653 37995
rect 6687 37992 6699 37995
rect 6687 37964 6914 37992
rect 6687 37961 6699 37964
rect 6641 37955 6699 37961
rect 6886 37924 6914 37964
rect 7009 37927 7067 37933
rect 7009 37924 7021 37927
rect 6886 37896 7021 37924
rect 7009 37893 7021 37896
rect 7055 37893 7067 37927
rect 7009 37887 7067 37893
rect 8018 37884 8024 37936
rect 8076 37884 8082 37936
rect 5307 37828 5488 37856
rect 5307 37825 5319 37828
rect 5261 37819 5319 37825
rect 6454 37816 6460 37868
rect 6512 37816 6518 37868
rect 5902 37748 5908 37800
rect 5960 37748 5966 37800
rect 6086 37748 6092 37800
rect 6144 37748 6150 37800
rect 6730 37748 6736 37800
rect 6788 37748 6794 37800
rect 7098 37612 7104 37664
rect 7156 37652 7162 37664
rect 7742 37652 7748 37664
rect 7156 37624 7748 37652
rect 7156 37612 7162 37624
rect 7742 37612 7748 37624
rect 7800 37652 7806 37664
rect 8481 37655 8539 37661
rect 8481 37652 8493 37655
rect 7800 37624 8493 37652
rect 7800 37612 7806 37624
rect 8481 37621 8493 37624
rect 8527 37621 8539 37655
rect 8481 37615 8539 37621
rect 1104 37562 8832 37584
rect 1104 37510 2350 37562
rect 2402 37510 2414 37562
rect 2466 37510 2478 37562
rect 2530 37510 2542 37562
rect 2594 37510 2606 37562
rect 2658 37510 7350 37562
rect 7402 37510 7414 37562
rect 7466 37510 7478 37562
rect 7530 37510 7542 37562
rect 7594 37510 7606 37562
rect 7658 37510 8832 37562
rect 1104 37488 8832 37510
rect 6454 37408 6460 37460
rect 6512 37448 6518 37460
rect 6733 37451 6791 37457
rect 6733 37448 6745 37451
rect 6512 37420 6745 37448
rect 6512 37408 6518 37420
rect 6733 37417 6745 37420
rect 6779 37417 6791 37451
rect 6733 37411 6791 37417
rect 5997 37315 6055 37321
rect 5997 37281 6009 37315
rect 6043 37312 6055 37315
rect 6086 37312 6092 37324
rect 6043 37284 6092 37312
rect 6043 37281 6055 37284
rect 5997 37275 6055 37281
rect 6086 37272 6092 37284
rect 6144 37272 6150 37324
rect 7190 37272 7196 37324
rect 7248 37312 7254 37324
rect 7285 37315 7343 37321
rect 7285 37312 7297 37315
rect 7248 37284 7297 37312
rect 7248 37272 7254 37284
rect 7285 37281 7297 37284
rect 7331 37281 7343 37315
rect 7285 37275 7343 37281
rect 5261 37247 5319 37253
rect 5261 37213 5273 37247
rect 5307 37244 5319 37247
rect 5307 37216 5396 37244
rect 5307 37213 5319 37216
rect 5261 37207 5319 37213
rect 5074 37068 5080 37120
rect 5132 37068 5138 37120
rect 5368 37117 5396 37216
rect 7098 37204 7104 37256
rect 7156 37204 7162 37256
rect 5721 37179 5779 37185
rect 5721 37145 5733 37179
rect 5767 37176 5779 37179
rect 5902 37176 5908 37188
rect 5767 37148 5908 37176
rect 5767 37145 5779 37148
rect 5721 37139 5779 37145
rect 5902 37136 5908 37148
rect 5960 37176 5966 37188
rect 7193 37179 7251 37185
rect 7193 37176 7205 37179
rect 5960 37148 7205 37176
rect 5960 37136 5966 37148
rect 7193 37145 7205 37148
rect 7239 37145 7251 37179
rect 7193 37139 7251 37145
rect 5353 37111 5411 37117
rect 5353 37077 5365 37111
rect 5399 37077 5411 37111
rect 5353 37071 5411 37077
rect 5813 37111 5871 37117
rect 5813 37077 5825 37111
rect 5859 37108 5871 37111
rect 6178 37108 6184 37120
rect 5859 37080 6184 37108
rect 5859 37077 5871 37080
rect 5813 37071 5871 37077
rect 6178 37068 6184 37080
rect 6236 37068 6242 37120
rect 1104 37018 8832 37040
rect 1104 36966 3010 37018
rect 3062 36966 3074 37018
rect 3126 36966 3138 37018
rect 3190 36966 3202 37018
rect 3254 36966 3266 37018
rect 3318 36966 8010 37018
rect 8062 36966 8074 37018
rect 8126 36966 8138 37018
rect 8190 36966 8202 37018
rect 8254 36966 8266 37018
rect 8318 36966 8832 37018
rect 1104 36944 8832 36966
rect 5074 36864 5080 36916
rect 5132 36864 5138 36916
rect 6178 36864 6184 36916
rect 6236 36864 6242 36916
rect 6641 36907 6699 36913
rect 6641 36873 6653 36907
rect 6687 36904 6699 36907
rect 6687 36876 6914 36904
rect 6687 36873 6699 36876
rect 6641 36867 6699 36873
rect 4709 36839 4767 36845
rect 4709 36805 4721 36839
rect 4755 36836 4767 36839
rect 5092 36836 5120 36864
rect 4755 36808 5120 36836
rect 6886 36836 6914 36876
rect 7926 36864 7932 36916
rect 7984 36904 7990 36916
rect 7984 36876 8156 36904
rect 7984 36864 7990 36876
rect 7009 36839 7067 36845
rect 7009 36836 7021 36839
rect 6886 36808 7021 36836
rect 4755 36805 4767 36808
rect 4709 36799 4767 36805
rect 7009 36805 7021 36808
rect 7055 36805 7067 36839
rect 7009 36799 7067 36805
rect 4430 36660 4436 36712
rect 4488 36660 4494 36712
rect 5828 36632 5856 36754
rect 6454 36728 6460 36780
rect 6512 36728 6518 36780
rect 6730 36660 6736 36712
rect 6788 36660 6794 36712
rect 7742 36700 7748 36712
rect 6840 36672 7748 36700
rect 5994 36632 6000 36644
rect 5828 36604 6000 36632
rect 5994 36592 6000 36604
rect 6052 36632 6058 36644
rect 6840 36632 6868 36672
rect 7742 36660 7748 36672
rect 7800 36700 7806 36712
rect 8128 36700 8156 36876
rect 7800 36672 8156 36700
rect 7800 36660 7806 36672
rect 6052 36604 6868 36632
rect 6052 36592 6058 36604
rect 8481 36567 8539 36573
rect 8481 36533 8493 36567
rect 8527 36564 8539 36567
rect 8527 36536 8892 36564
rect 8527 36533 8539 36536
rect 8481 36527 8539 36533
rect 1104 36474 8832 36496
rect 1104 36422 2350 36474
rect 2402 36422 2414 36474
rect 2466 36422 2478 36474
rect 2530 36422 2542 36474
rect 2594 36422 2606 36474
rect 2658 36422 7350 36474
rect 7402 36422 7414 36474
rect 7466 36422 7478 36474
rect 7530 36422 7542 36474
rect 7594 36422 7606 36474
rect 7658 36422 8832 36474
rect 1104 36400 8832 36422
rect 6454 36320 6460 36372
rect 6512 36360 6518 36372
rect 6641 36363 6699 36369
rect 6641 36360 6653 36363
rect 6512 36332 6653 36360
rect 6512 36320 6518 36332
rect 6641 36329 6653 36332
rect 6687 36329 6699 36363
rect 6641 36323 6699 36329
rect 8386 36320 8392 36372
rect 8444 36320 8450 36372
rect 6178 36184 6184 36236
rect 6236 36224 6242 36236
rect 7101 36227 7159 36233
rect 7101 36224 7113 36227
rect 6236 36196 7113 36224
rect 6236 36184 6242 36196
rect 7101 36193 7113 36196
rect 7147 36193 7159 36227
rect 7101 36187 7159 36193
rect 7190 36184 7196 36236
rect 7248 36184 7254 36236
rect 7009 36159 7067 36165
rect 7009 36125 7021 36159
rect 7055 36156 7067 36159
rect 8205 36159 8263 36165
rect 8205 36156 8217 36159
rect 7055 36128 8217 36156
rect 7055 36125 7067 36128
rect 7009 36119 7067 36125
rect 8205 36125 8217 36128
rect 8251 36156 8263 36159
rect 8864 36156 8892 36536
rect 8251 36128 8892 36156
rect 8251 36125 8263 36128
rect 8205 36119 8263 36125
rect 1104 35930 8832 35952
rect 1104 35878 3010 35930
rect 3062 35878 3074 35930
rect 3126 35878 3138 35930
rect 3190 35878 3202 35930
rect 3254 35878 3266 35930
rect 3318 35878 8010 35930
rect 8062 35878 8074 35930
rect 8126 35878 8138 35930
rect 8190 35878 8202 35930
rect 8254 35878 8266 35930
rect 8318 35878 8832 35930
rect 1104 35856 8832 35878
rect 5813 35819 5871 35825
rect 5813 35785 5825 35819
rect 5859 35816 5871 35819
rect 6178 35816 6184 35828
rect 5859 35788 6184 35816
rect 5859 35785 5871 35788
rect 5813 35779 5871 35785
rect 6178 35776 6184 35788
rect 6236 35776 6242 35828
rect 5261 35683 5319 35689
rect 5261 35649 5273 35683
rect 5307 35680 5319 35683
rect 5307 35652 5488 35680
rect 5307 35649 5319 35652
rect 5261 35643 5319 35649
rect 5460 35553 5488 35652
rect 8018 35640 8024 35692
rect 8076 35680 8082 35692
rect 8205 35683 8263 35689
rect 8205 35680 8217 35683
rect 8076 35652 8217 35680
rect 8076 35640 8082 35652
rect 8205 35649 8217 35652
rect 8251 35649 8263 35683
rect 8205 35643 8263 35649
rect 5902 35572 5908 35624
rect 5960 35572 5966 35624
rect 6086 35572 6092 35624
rect 6144 35572 6150 35624
rect 5445 35547 5503 35553
rect 5445 35513 5457 35547
rect 5491 35513 5503 35547
rect 5445 35507 5503 35513
rect 4982 35436 4988 35488
rect 5040 35476 5046 35488
rect 5077 35479 5135 35485
rect 5077 35476 5089 35479
rect 5040 35448 5089 35476
rect 5040 35436 5046 35448
rect 5077 35445 5089 35448
rect 5123 35445 5135 35479
rect 5077 35439 5135 35445
rect 8386 35436 8392 35488
rect 8444 35436 8450 35488
rect 1104 35386 8832 35408
rect 1104 35334 2350 35386
rect 2402 35334 2414 35386
rect 2466 35334 2478 35386
rect 2530 35334 2542 35386
rect 2594 35334 2606 35386
rect 2658 35334 7350 35386
rect 7402 35334 7414 35386
rect 7466 35334 7478 35386
rect 7530 35334 7542 35386
rect 7594 35334 7606 35386
rect 7658 35334 8832 35386
rect 1104 35312 8832 35334
rect 5902 35232 5908 35284
rect 5960 35272 5966 35284
rect 6365 35275 6423 35281
rect 6365 35272 6377 35275
rect 5960 35244 6377 35272
rect 5960 35232 5966 35244
rect 6365 35241 6377 35244
rect 6411 35241 6423 35275
rect 6365 35235 6423 35241
rect 4893 35139 4951 35145
rect 4893 35105 4905 35139
rect 4939 35136 4951 35139
rect 4982 35136 4988 35148
rect 4939 35108 4988 35136
rect 4939 35105 4951 35108
rect 4893 35099 4951 35105
rect 4982 35096 4988 35108
rect 5040 35096 5046 35148
rect 4430 35028 4436 35080
rect 4488 35068 4494 35080
rect 4617 35071 4675 35077
rect 4617 35068 4629 35071
rect 4488 35040 4629 35068
rect 4488 35028 4494 35040
rect 4617 35037 4629 35040
rect 4663 35037 4675 35071
rect 4617 35031 4675 35037
rect 4632 35000 4660 35031
rect 6454 35028 6460 35080
rect 6512 35028 6518 35080
rect 6730 35028 6736 35080
rect 6788 35028 6794 35080
rect 6178 35000 6184 35012
rect 4632 34972 4844 35000
rect 6118 34972 6184 35000
rect 4816 34944 4844 34972
rect 6178 34960 6184 34972
rect 6236 34960 6242 35012
rect 7009 35003 7067 35009
rect 7009 35000 7021 35003
rect 6886 34972 7021 35000
rect 4798 34892 4804 34944
rect 4856 34892 4862 34944
rect 6641 34935 6699 34941
rect 6641 34901 6653 34935
rect 6687 34932 6699 34935
rect 6886 34932 6914 34972
rect 7009 34969 7021 34972
rect 7055 34969 7067 35003
rect 7009 34963 7067 34969
rect 7282 34960 7288 35012
rect 7340 35000 7346 35012
rect 7340 34972 7498 35000
rect 7340 34960 7346 34972
rect 6687 34904 6914 34932
rect 6687 34901 6699 34904
rect 6641 34895 6699 34901
rect 7098 34892 7104 34944
rect 7156 34932 7162 34944
rect 8018 34932 8024 34944
rect 7156 34904 8024 34932
rect 7156 34892 7162 34904
rect 8018 34892 8024 34904
rect 8076 34932 8082 34944
rect 8481 34935 8539 34941
rect 8481 34932 8493 34935
rect 8076 34904 8493 34932
rect 8076 34892 8082 34904
rect 8481 34901 8493 34904
rect 8527 34901 8539 34935
rect 8481 34895 8539 34901
rect 1104 34842 8832 34864
rect 1104 34790 3010 34842
rect 3062 34790 3074 34842
rect 3126 34790 3138 34842
rect 3190 34790 3202 34842
rect 3254 34790 3266 34842
rect 3318 34790 8010 34842
rect 8062 34790 8074 34842
rect 8126 34790 8138 34842
rect 8190 34790 8202 34842
rect 8254 34790 8266 34842
rect 8318 34790 8832 34842
rect 1104 34768 8832 34790
rect 4617 34663 4675 34669
rect 4617 34629 4629 34663
rect 4663 34660 4675 34663
rect 4663 34632 6868 34660
rect 4663 34629 4675 34632
rect 4617 34623 4675 34629
rect 6840 34604 6868 34632
rect 5442 34552 5448 34604
rect 5500 34592 5506 34604
rect 5813 34595 5871 34601
rect 5813 34592 5825 34595
rect 5500 34564 5825 34592
rect 5500 34552 5506 34564
rect 5813 34561 5825 34564
rect 5859 34561 5871 34595
rect 5813 34555 5871 34561
rect 6822 34552 6828 34604
rect 6880 34552 6886 34604
rect 4798 34484 4804 34536
rect 4856 34524 4862 34536
rect 5353 34527 5411 34533
rect 5353 34524 5365 34527
rect 4856 34496 5365 34524
rect 4856 34484 4862 34496
rect 5353 34493 5365 34496
rect 5399 34493 5411 34527
rect 5353 34487 5411 34493
rect 6730 34484 6736 34536
rect 6788 34524 6794 34536
rect 7561 34527 7619 34533
rect 7561 34524 7573 34527
rect 6788 34496 7573 34524
rect 6788 34484 6794 34496
rect 7561 34493 7573 34496
rect 7607 34493 7619 34527
rect 7561 34487 7619 34493
rect 5626 34348 5632 34400
rect 5684 34348 5690 34400
rect 1104 34298 8832 34320
rect 1104 34246 2350 34298
rect 2402 34246 2414 34298
rect 2466 34246 2478 34298
rect 2530 34246 2542 34298
rect 2594 34246 2606 34298
rect 2658 34246 7350 34298
rect 7402 34246 7414 34298
rect 7466 34246 7478 34298
rect 7530 34246 7542 34298
rect 7594 34246 7606 34298
rect 7658 34246 8832 34298
rect 1104 34224 8832 34246
rect 5064 34187 5122 34193
rect 5064 34153 5076 34187
rect 5110 34184 5122 34187
rect 5626 34184 5632 34196
rect 5110 34156 5632 34184
rect 5110 34153 5122 34156
rect 5064 34147 5122 34153
rect 5626 34144 5632 34156
rect 5684 34144 5690 34196
rect 4798 34076 4804 34128
rect 4856 34076 4862 34128
rect 4816 34048 4844 34076
rect 6733 34051 6791 34057
rect 6733 34048 6745 34051
rect 4816 34020 6745 34048
rect 6733 34017 6745 34020
rect 6779 34017 6791 34051
rect 6733 34011 6791 34017
rect 7006 34008 7012 34060
rect 7064 34048 7070 34060
rect 7374 34048 7380 34060
rect 7064 34020 7380 34048
rect 7064 34008 7070 34020
rect 7374 34008 7380 34020
rect 7432 34008 7438 34060
rect 4801 33983 4859 33989
rect 4801 33949 4813 33983
rect 4847 33949 4859 33983
rect 4801 33943 4859 33949
rect 4816 33844 4844 33943
rect 6178 33940 6184 33992
rect 6236 33980 6242 33992
rect 6236 33952 6776 33980
rect 6236 33940 6242 33952
rect 6748 33912 6776 33952
rect 6380 33884 6684 33912
rect 6748 33884 6914 33912
rect 6380 33844 6408 33884
rect 4816 33816 6408 33844
rect 6546 33804 6552 33856
rect 6604 33804 6610 33856
rect 6656 33844 6684 33884
rect 6730 33844 6736 33856
rect 6656 33816 6736 33844
rect 6730 33804 6736 33816
rect 6788 33804 6794 33856
rect 6886 33844 6914 33884
rect 7006 33872 7012 33924
rect 7064 33872 7070 33924
rect 7208 33884 7498 33912
rect 7208 33856 7236 33884
rect 7190 33844 7196 33856
rect 6886 33816 7196 33844
rect 7190 33804 7196 33816
rect 7248 33804 7254 33856
rect 7926 33804 7932 33856
rect 7984 33844 7990 33856
rect 8481 33847 8539 33853
rect 8481 33844 8493 33847
rect 7984 33816 8493 33844
rect 7984 33804 7990 33816
rect 8481 33813 8493 33816
rect 8527 33813 8539 33847
rect 8481 33807 8539 33813
rect 1104 33754 8832 33776
rect 1104 33702 3010 33754
rect 3062 33702 3074 33754
rect 3126 33702 3138 33754
rect 3190 33702 3202 33754
rect 3254 33702 3266 33754
rect 3318 33702 8010 33754
rect 8062 33702 8074 33754
rect 8126 33702 8138 33754
rect 8190 33702 8202 33754
rect 8254 33702 8266 33754
rect 8318 33702 8832 33754
rect 1104 33680 8832 33702
rect 5442 33600 5448 33652
rect 5500 33600 5506 33652
rect 5810 33600 5816 33652
rect 5868 33600 5874 33652
rect 6454 33600 6460 33652
rect 6512 33640 6518 33652
rect 6733 33643 6791 33649
rect 6733 33640 6745 33643
rect 6512 33612 6745 33640
rect 6512 33600 6518 33612
rect 6733 33609 6745 33612
rect 6779 33609 6791 33643
rect 6733 33603 6791 33609
rect 7098 33600 7104 33652
rect 7156 33600 7162 33652
rect 7926 33600 7932 33652
rect 7984 33600 7990 33652
rect 5828 33504 5856 33600
rect 5905 33575 5963 33581
rect 5905 33541 5917 33575
rect 5951 33572 5963 33575
rect 6546 33572 6552 33584
rect 5951 33544 6552 33572
rect 5951 33541 5963 33544
rect 5905 33535 5963 33541
rect 6546 33532 6552 33544
rect 6604 33572 6610 33584
rect 8021 33575 8079 33581
rect 8021 33572 8033 33575
rect 6604 33544 8033 33572
rect 6604 33532 6610 33544
rect 8021 33541 8033 33544
rect 8067 33541 8079 33575
rect 8021 33535 8079 33541
rect 7193 33507 7251 33513
rect 5828 33476 6914 33504
rect 6086 33396 6092 33448
rect 6144 33396 6150 33448
rect 6886 33436 6914 33476
rect 7193 33473 7205 33507
rect 7239 33473 7251 33507
rect 7193 33467 7251 33473
rect 7208 33436 7236 33467
rect 6886 33408 7236 33436
rect 7374 33396 7380 33448
rect 7432 33436 7438 33448
rect 8018 33436 8024 33448
rect 7432 33408 8024 33436
rect 7432 33396 7438 33408
rect 8018 33396 8024 33408
rect 8076 33436 8082 33448
rect 8113 33439 8171 33445
rect 8113 33436 8125 33439
rect 8076 33408 8125 33436
rect 8076 33396 8082 33408
rect 8113 33405 8125 33408
rect 8159 33405 8171 33439
rect 8113 33399 8171 33405
rect 7190 33260 7196 33312
rect 7248 33300 7254 33312
rect 7561 33303 7619 33309
rect 7561 33300 7573 33303
rect 7248 33272 7573 33300
rect 7248 33260 7254 33272
rect 7561 33269 7573 33272
rect 7607 33269 7619 33303
rect 7561 33263 7619 33269
rect 1104 33210 8832 33232
rect 1104 33158 2350 33210
rect 2402 33158 2414 33210
rect 2466 33158 2478 33210
rect 2530 33158 2542 33210
rect 2594 33158 2606 33210
rect 2658 33158 7350 33210
rect 7402 33158 7414 33210
rect 7466 33158 7478 33210
rect 7530 33158 7542 33210
rect 7594 33158 7606 33210
rect 7658 33158 8832 33210
rect 1104 33136 8832 33158
rect 7006 33056 7012 33108
rect 7064 33056 7070 33108
rect 7561 33099 7619 33105
rect 7561 33065 7573 33099
rect 7607 33096 7619 33099
rect 7742 33096 7748 33108
rect 7607 33068 7748 33096
rect 7607 33065 7619 33068
rect 7561 33059 7619 33065
rect 7742 33056 7748 33068
rect 7800 33056 7806 33108
rect 7926 33056 7932 33108
rect 7984 33056 7990 33108
rect 7190 32852 7196 32904
rect 7248 32852 7254 32904
rect 7653 32895 7711 32901
rect 7653 32861 7665 32895
rect 7699 32892 7711 32895
rect 7944 32892 7972 33056
rect 7699 32864 7972 32892
rect 7699 32861 7711 32864
rect 7653 32855 7711 32861
rect 7742 32784 7748 32836
rect 7800 32824 7806 32836
rect 7929 32827 7987 32833
rect 7929 32824 7941 32827
rect 7800 32796 7941 32824
rect 7800 32784 7806 32796
rect 7929 32793 7941 32796
rect 7975 32793 7987 32827
rect 7929 32787 7987 32793
rect 8205 32759 8263 32765
rect 8205 32725 8217 32759
rect 8251 32756 8263 32759
rect 8662 32756 8668 32768
rect 8251 32728 8668 32756
rect 8251 32725 8263 32728
rect 8205 32719 8263 32725
rect 8662 32716 8668 32728
rect 8720 32716 8726 32768
rect 1104 32666 8832 32688
rect 1104 32614 3010 32666
rect 3062 32614 3074 32666
rect 3126 32614 3138 32666
rect 3190 32614 3202 32666
rect 3254 32614 3266 32666
rect 3318 32614 8010 32666
rect 8062 32614 8074 32666
rect 8126 32614 8138 32666
rect 8190 32614 8202 32666
rect 8254 32614 8266 32666
rect 8318 32614 8832 32666
rect 1104 32592 8832 32614
rect 6641 32555 6699 32561
rect 6641 32521 6653 32555
rect 6687 32552 6699 32555
rect 6687 32524 6914 32552
rect 6687 32521 6699 32524
rect 6641 32515 6699 32521
rect 6886 32484 6914 32524
rect 7009 32487 7067 32493
rect 7009 32484 7021 32487
rect 5934 32456 6592 32484
rect 6886 32456 7021 32484
rect 6564 32428 6592 32456
rect 7009 32453 7021 32456
rect 7055 32453 7067 32487
rect 7009 32447 7067 32453
rect 7098 32444 7104 32496
rect 7156 32484 7162 32496
rect 7156 32456 7498 32484
rect 7156 32444 7162 32456
rect 6454 32376 6460 32428
rect 6512 32376 6518 32428
rect 6546 32376 6552 32428
rect 6604 32376 6610 32428
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32317 4491 32351
rect 4433 32311 4491 32317
rect 4448 32212 4476 32311
rect 4706 32308 4712 32360
rect 4764 32308 4770 32360
rect 6730 32308 6736 32360
rect 6788 32308 6794 32360
rect 4798 32212 4804 32224
rect 4448 32184 4804 32212
rect 4798 32172 4804 32184
rect 4856 32172 4862 32224
rect 6178 32172 6184 32224
rect 6236 32172 6242 32224
rect 7098 32172 7104 32224
rect 7156 32212 7162 32224
rect 7742 32212 7748 32224
rect 7156 32184 7748 32212
rect 7156 32172 7162 32184
rect 7742 32172 7748 32184
rect 7800 32212 7806 32224
rect 8481 32215 8539 32221
rect 8481 32212 8493 32215
rect 7800 32184 8493 32212
rect 7800 32172 7806 32184
rect 8481 32181 8493 32184
rect 8527 32181 8539 32215
rect 8481 32175 8539 32181
rect 1104 32122 8832 32144
rect 1104 32070 2350 32122
rect 2402 32070 2414 32122
rect 2466 32070 2478 32122
rect 2530 32070 2542 32122
rect 2594 32070 2606 32122
rect 2658 32070 7350 32122
rect 7402 32070 7414 32122
rect 7466 32070 7478 32122
rect 7530 32070 7542 32122
rect 7594 32070 7606 32122
rect 7658 32070 8832 32122
rect 1104 32048 8832 32070
rect 4706 31968 4712 32020
rect 4764 32008 4770 32020
rect 5077 32011 5135 32017
rect 5077 32008 5089 32011
rect 4764 31980 5089 32008
rect 4764 31968 4770 31980
rect 5077 31977 5089 31980
rect 5123 31977 5135 32011
rect 5077 31971 5135 31977
rect 6454 31968 6460 32020
rect 6512 32008 6518 32020
rect 6733 32011 6791 32017
rect 6733 32008 6745 32011
rect 6512 31980 6745 32008
rect 6512 31968 6518 31980
rect 6733 31977 6745 31980
rect 6779 31977 6791 32011
rect 6733 31971 6791 31977
rect 5537 31943 5595 31949
rect 5537 31909 5549 31943
rect 5583 31909 5595 31943
rect 5537 31903 5595 31909
rect 5261 31807 5319 31813
rect 5261 31773 5273 31807
rect 5307 31804 5319 31807
rect 5552 31804 5580 31903
rect 5994 31832 6000 31884
rect 6052 31872 6058 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 6052 31844 6101 31872
rect 6052 31832 6058 31844
rect 6089 31841 6101 31844
rect 6135 31841 6147 31875
rect 7193 31875 7251 31881
rect 7193 31872 7205 31875
rect 6089 31835 6147 31841
rect 6932 31844 7205 31872
rect 6932 31816 6960 31844
rect 7193 31841 7205 31844
rect 7239 31841 7251 31875
rect 7193 31835 7251 31841
rect 7377 31875 7435 31881
rect 7377 31841 7389 31875
rect 7423 31872 7435 31875
rect 7742 31872 7748 31884
rect 7423 31844 7748 31872
rect 7423 31841 7435 31844
rect 7377 31835 7435 31841
rect 7742 31832 7748 31844
rect 7800 31872 7806 31884
rect 7926 31872 7932 31884
rect 7800 31844 7932 31872
rect 7800 31832 7806 31844
rect 7926 31832 7932 31844
rect 7984 31832 7990 31884
rect 6914 31804 6920 31816
rect 5307 31776 5580 31804
rect 5307 31773 5319 31776
rect 5261 31767 5319 31773
rect 6886 31764 6920 31804
rect 6972 31764 6978 31816
rect 7098 31764 7104 31816
rect 7156 31764 7162 31816
rect 5445 31739 5503 31745
rect 5445 31705 5457 31739
rect 5491 31736 5503 31739
rect 5905 31739 5963 31745
rect 5905 31736 5917 31739
rect 5491 31708 5917 31736
rect 5491 31705 5503 31708
rect 5445 31699 5503 31705
rect 5905 31705 5917 31708
rect 5951 31736 5963 31739
rect 6886 31736 6914 31764
rect 5951 31708 6914 31736
rect 5951 31705 5963 31708
rect 5905 31699 5963 31705
rect 5997 31671 6055 31677
rect 5997 31637 6009 31671
rect 6043 31668 6055 31671
rect 6178 31668 6184 31680
rect 6043 31640 6184 31668
rect 6043 31637 6055 31640
rect 5997 31631 6055 31637
rect 6178 31628 6184 31640
rect 6236 31628 6242 31680
rect 1104 31578 8832 31600
rect 1104 31526 3010 31578
rect 3062 31526 3074 31578
rect 3126 31526 3138 31578
rect 3190 31526 3202 31578
rect 3254 31526 3266 31578
rect 3318 31526 8010 31578
rect 8062 31526 8074 31578
rect 8126 31526 8138 31578
rect 8190 31526 8202 31578
rect 8254 31526 8266 31578
rect 8318 31526 8832 31578
rect 1104 31504 8832 31526
rect 6641 31467 6699 31473
rect 6641 31433 6653 31467
rect 6687 31433 6699 31467
rect 6641 31427 6699 31433
rect 6656 31396 6684 31427
rect 7009 31399 7067 31405
rect 7009 31396 7021 31399
rect 6656 31368 7021 31396
rect 7009 31365 7021 31368
rect 7055 31365 7067 31399
rect 7009 31359 7067 31365
rect 8018 31356 8024 31408
rect 8076 31356 8082 31408
rect 6454 31288 6460 31340
rect 6512 31288 6518 31340
rect 6730 31220 6736 31272
rect 6788 31220 6794 31272
rect 8481 31127 8539 31133
rect 8481 31093 8493 31127
rect 8527 31124 8539 31127
rect 8527 31096 8892 31124
rect 8527 31093 8539 31096
rect 8481 31087 8539 31093
rect 1104 31034 8832 31056
rect 1104 30982 2350 31034
rect 2402 30982 2414 31034
rect 2466 30982 2478 31034
rect 2530 30982 2542 31034
rect 2594 30982 2606 31034
rect 2658 30982 7350 31034
rect 7402 30982 7414 31034
rect 7466 30982 7478 31034
rect 7530 30982 7542 31034
rect 7594 30982 7606 31034
rect 7658 30982 8832 31034
rect 1104 30960 8832 30982
rect 6454 30880 6460 30932
rect 6512 30920 6518 30932
rect 6733 30923 6791 30929
rect 6733 30920 6745 30923
rect 6512 30892 6745 30920
rect 6512 30880 6518 30892
rect 6733 30889 6745 30892
rect 6779 30889 6791 30923
rect 6733 30883 6791 30889
rect 7929 30923 7987 30929
rect 7929 30889 7941 30923
rect 7975 30920 7987 30923
rect 8018 30920 8024 30932
rect 7975 30892 8024 30920
rect 7975 30889 7987 30892
rect 7929 30883 7987 30889
rect 7944 30852 7972 30883
rect 8018 30880 8024 30892
rect 8076 30880 8082 30932
rect 8386 30880 8392 30932
rect 8444 30880 8450 30932
rect 6380 30824 7972 30852
rect 4798 30744 4804 30796
rect 4856 30744 4862 30796
rect 6380 30716 6408 30824
rect 6454 30744 6460 30796
rect 6512 30784 6518 30796
rect 7193 30787 7251 30793
rect 7193 30784 7205 30787
rect 6512 30756 7205 30784
rect 6512 30744 6518 30756
rect 7193 30753 7205 30756
rect 7239 30753 7251 30787
rect 7193 30747 7251 30753
rect 7377 30787 7435 30793
rect 7377 30753 7389 30787
rect 7423 30784 7435 30787
rect 7742 30784 7748 30796
rect 7423 30756 7748 30784
rect 7423 30753 7435 30756
rect 7377 30747 7435 30753
rect 7742 30744 7748 30756
rect 7800 30744 7806 30796
rect 6210 30688 6408 30716
rect 6546 30676 6552 30728
rect 6604 30676 6610 30728
rect 7101 30719 7159 30725
rect 7101 30685 7113 30719
rect 7147 30716 7159 30719
rect 8205 30719 8263 30725
rect 8205 30716 8217 30719
rect 7147 30688 8217 30716
rect 7147 30685 7159 30688
rect 7101 30679 7159 30685
rect 8205 30685 8217 30688
rect 8251 30716 8263 30719
rect 8864 30716 8892 31096
rect 8251 30688 8892 30716
rect 8251 30685 8263 30688
rect 8205 30679 8263 30685
rect 5074 30608 5080 30660
rect 5132 30608 5138 30660
rect 6564 30648 6592 30676
rect 7653 30651 7711 30657
rect 7653 30648 7665 30651
rect 6564 30620 7665 30648
rect 7653 30617 7665 30620
rect 7699 30617 7711 30651
rect 7653 30611 7711 30617
rect 6549 30583 6607 30589
rect 6549 30549 6561 30583
rect 6595 30580 6607 30583
rect 6638 30580 6644 30592
rect 6595 30552 6644 30580
rect 6595 30549 6607 30552
rect 6549 30543 6607 30549
rect 6638 30540 6644 30552
rect 6696 30540 6702 30592
rect 1104 30490 8832 30512
rect 1104 30438 3010 30490
rect 3062 30438 3074 30490
rect 3126 30438 3138 30490
rect 3190 30438 3202 30490
rect 3254 30438 3266 30490
rect 3318 30438 8010 30490
rect 8062 30438 8074 30490
rect 8126 30438 8138 30490
rect 8190 30438 8202 30490
rect 8254 30438 8266 30490
rect 8318 30438 8832 30490
rect 1104 30416 8832 30438
rect 5074 30336 5080 30388
rect 5132 30376 5138 30388
rect 5169 30379 5227 30385
rect 5169 30376 5181 30379
rect 5132 30348 5181 30376
rect 5132 30336 5138 30348
rect 5169 30345 5181 30348
rect 5215 30345 5227 30379
rect 5169 30339 5227 30345
rect 6178 30336 6184 30388
rect 6236 30376 6242 30388
rect 6454 30376 6460 30388
rect 6236 30348 6460 30376
rect 6236 30336 6242 30348
rect 6454 30336 6460 30348
rect 6512 30376 6518 30388
rect 6512 30348 6776 30376
rect 6512 30336 6518 30348
rect 6086 30268 6092 30320
rect 6144 30308 6150 30320
rect 6748 30317 6776 30348
rect 6733 30311 6791 30317
rect 6144 30280 6684 30308
rect 6144 30268 6150 30280
rect 5353 30243 5411 30249
rect 5353 30209 5365 30243
rect 5399 30240 5411 30243
rect 6656 30240 6684 30280
rect 6733 30277 6745 30311
rect 6779 30277 6791 30311
rect 6733 30271 6791 30277
rect 8205 30243 8263 30249
rect 5399 30212 6408 30240
rect 6656 30212 6960 30240
rect 5399 30209 5411 30212
rect 5353 30203 5411 30209
rect 6380 30113 6408 30212
rect 6638 30132 6644 30184
rect 6696 30172 6702 30184
rect 6932 30181 6960 30212
rect 8205 30209 8217 30243
rect 8251 30240 8263 30243
rect 8251 30212 8892 30240
rect 8251 30209 8263 30212
rect 8205 30203 8263 30209
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 6696 30144 6837 30172
rect 6696 30132 6702 30144
rect 6825 30141 6837 30144
rect 6871 30141 6883 30175
rect 6825 30135 6883 30141
rect 6917 30175 6975 30181
rect 6917 30141 6929 30175
rect 6963 30141 6975 30175
rect 6917 30135 6975 30141
rect 6365 30107 6423 30113
rect 6365 30073 6377 30107
rect 6411 30073 6423 30107
rect 6365 30067 6423 30073
rect 8386 29996 8392 30048
rect 8444 29996 8450 30048
rect 1104 29946 8832 29968
rect 1104 29894 2350 29946
rect 2402 29894 2414 29946
rect 2466 29894 2478 29946
rect 2530 29894 2542 29946
rect 2594 29894 2606 29946
rect 2658 29894 7350 29946
rect 7402 29894 7414 29946
rect 7466 29894 7478 29946
rect 7530 29894 7542 29946
rect 7594 29894 7606 29946
rect 7658 29894 8832 29946
rect 1104 29872 8832 29894
rect 6086 29656 6092 29708
rect 6144 29656 6150 29708
rect 6270 29656 6276 29708
rect 6328 29656 6334 29708
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29628 6055 29631
rect 6288 29628 6316 29656
rect 6043 29600 6316 29628
rect 6043 29597 6055 29600
rect 5997 29591 6055 29597
rect 6454 29588 6460 29640
rect 6512 29588 6518 29640
rect 6730 29588 6736 29640
rect 6788 29588 6794 29640
rect 8018 29588 8024 29640
rect 8076 29628 8082 29640
rect 8076 29600 8142 29628
rect 8076 29588 8082 29600
rect 7009 29563 7067 29569
rect 7009 29560 7021 29563
rect 6656 29532 7021 29560
rect 5258 29452 5264 29504
rect 5316 29492 5322 29504
rect 5537 29495 5595 29501
rect 5537 29492 5549 29495
rect 5316 29464 5549 29492
rect 5316 29452 5322 29464
rect 5537 29461 5549 29464
rect 5583 29461 5595 29495
rect 5537 29455 5595 29461
rect 5902 29452 5908 29504
rect 5960 29452 5966 29504
rect 6656 29501 6684 29532
rect 7009 29529 7021 29532
rect 7055 29529 7067 29563
rect 7009 29523 7067 29529
rect 6641 29495 6699 29501
rect 6641 29461 6653 29495
rect 6687 29461 6699 29495
rect 6641 29455 6699 29461
rect 8481 29495 8539 29501
rect 8481 29461 8493 29495
rect 8527 29492 8539 29495
rect 8864 29492 8892 30212
rect 8527 29464 8892 29492
rect 8527 29461 8539 29464
rect 8481 29455 8539 29461
rect 1104 29402 8832 29424
rect 1104 29350 3010 29402
rect 3062 29350 3074 29402
rect 3126 29350 3138 29402
rect 3190 29350 3202 29402
rect 3254 29350 3266 29402
rect 3318 29350 8010 29402
rect 8062 29350 8074 29402
rect 8126 29350 8138 29402
rect 8190 29350 8202 29402
rect 8254 29350 8266 29402
rect 8318 29350 8832 29402
rect 1104 29328 8832 29350
rect 5258 29248 5264 29300
rect 5316 29248 5322 29300
rect 5445 29291 5503 29297
rect 5445 29257 5457 29291
rect 5491 29257 5503 29291
rect 5445 29251 5503 29257
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29152 5135 29155
rect 5276 29152 5304 29248
rect 5123 29124 5304 29152
rect 5353 29155 5411 29161
rect 5123 29121 5135 29124
rect 5077 29115 5135 29121
rect 5353 29121 5365 29155
rect 5399 29152 5411 29155
rect 5460 29152 5488 29251
rect 6454 29248 6460 29300
rect 6512 29288 6518 29300
rect 6825 29291 6883 29297
rect 6825 29288 6837 29291
rect 6512 29260 6837 29288
rect 6512 29248 6518 29260
rect 6825 29257 6837 29260
rect 6871 29257 6883 29291
rect 6825 29251 6883 29257
rect 7193 29291 7251 29297
rect 7193 29257 7205 29291
rect 7239 29288 7251 29291
rect 8864 29288 8892 29464
rect 7239 29260 8892 29288
rect 7239 29257 7251 29260
rect 7193 29251 7251 29257
rect 5813 29223 5871 29229
rect 5813 29189 5825 29223
rect 5859 29220 5871 29223
rect 6638 29220 6644 29232
rect 5859 29192 6644 29220
rect 5859 29189 5871 29192
rect 5813 29183 5871 29189
rect 6638 29180 6644 29192
rect 6696 29220 6702 29232
rect 7285 29223 7343 29229
rect 7285 29220 7297 29223
rect 6696 29192 7297 29220
rect 6696 29180 6702 29192
rect 7285 29189 7297 29192
rect 7331 29189 7343 29223
rect 7285 29183 7343 29189
rect 5399 29124 5488 29152
rect 5399 29121 5411 29124
rect 5353 29115 5411 29121
rect 5902 29112 5908 29164
rect 5960 29152 5966 29164
rect 5960 29124 6592 29152
rect 5960 29112 5966 29124
rect 6564 29096 6592 29124
rect 6086 29044 6092 29096
rect 6144 29044 6150 29096
rect 6546 29044 6552 29096
rect 6604 29044 6610 29096
rect 7469 29087 7527 29093
rect 7469 29053 7481 29087
rect 7515 29084 7527 29087
rect 7742 29084 7748 29096
rect 7515 29056 7748 29084
rect 7515 29053 7527 29056
rect 7469 29047 7527 29053
rect 7190 28976 7196 29028
rect 7248 29016 7254 29028
rect 7484 29016 7512 29047
rect 7742 29044 7748 29056
rect 7800 29044 7806 29096
rect 7248 28988 7512 29016
rect 7248 28976 7254 28988
rect 4706 28908 4712 28960
rect 4764 28948 4770 28960
rect 4893 28951 4951 28957
rect 4893 28948 4905 28951
rect 4764 28920 4905 28948
rect 4764 28908 4770 28920
rect 4893 28917 4905 28920
rect 4939 28917 4951 28951
rect 4893 28911 4951 28917
rect 5166 28908 5172 28960
rect 5224 28908 5230 28960
rect 1104 28858 8832 28880
rect 1104 28806 2350 28858
rect 2402 28806 2414 28858
rect 2466 28806 2478 28858
rect 2530 28806 2542 28858
rect 2594 28806 2606 28858
rect 2658 28806 7350 28858
rect 7402 28806 7414 28858
rect 7466 28806 7478 28858
rect 7530 28806 7542 28858
rect 7594 28806 7606 28858
rect 7658 28806 8832 28858
rect 1104 28784 8832 28806
rect 4798 28568 4804 28620
rect 4856 28568 4862 28620
rect 5077 28611 5135 28617
rect 5077 28577 5089 28611
rect 5123 28608 5135 28611
rect 5166 28608 5172 28620
rect 5123 28580 5172 28608
rect 5123 28577 5135 28580
rect 5077 28571 5135 28577
rect 5166 28568 5172 28580
rect 5224 28568 5230 28620
rect 7098 28608 7104 28620
rect 6196 28580 7104 28608
rect 6086 28500 6092 28552
rect 6144 28540 6150 28552
rect 6196 28540 6224 28580
rect 7098 28568 7104 28580
rect 7156 28608 7162 28620
rect 7156 28580 8064 28608
rect 7156 28568 7162 28580
rect 8036 28552 8064 28580
rect 6144 28526 6224 28540
rect 6144 28512 6210 28526
rect 6144 28500 6150 28512
rect 6730 28500 6736 28552
rect 6788 28500 6794 28552
rect 8018 28500 8024 28552
rect 8076 28540 8082 28552
rect 8076 28512 8142 28540
rect 8076 28500 8082 28512
rect 7006 28432 7012 28484
rect 7064 28432 7070 28484
rect 6546 28364 6552 28416
rect 6604 28364 6610 28416
rect 8481 28407 8539 28413
rect 8481 28373 8493 28407
rect 8527 28404 8539 28407
rect 8527 28376 8892 28404
rect 8527 28373 8539 28376
rect 8481 28367 8539 28373
rect 1104 28314 8832 28336
rect 1104 28262 3010 28314
rect 3062 28262 3074 28314
rect 3126 28262 3138 28314
rect 3190 28262 3202 28314
rect 3254 28262 3266 28314
rect 3318 28262 8010 28314
rect 8062 28262 8074 28314
rect 8126 28262 8138 28314
rect 8190 28262 8202 28314
rect 8254 28262 8266 28314
rect 8318 28262 8832 28314
rect 1104 28240 8832 28262
rect 4798 28160 4804 28212
rect 4856 28160 4862 28212
rect 6086 28160 6092 28212
rect 6144 28160 6150 28212
rect 6181 28203 6239 28209
rect 6181 28169 6193 28203
rect 6227 28200 6239 28203
rect 6270 28200 6276 28212
rect 6227 28172 6276 28200
rect 6227 28169 6239 28172
rect 6181 28163 6239 28169
rect 6270 28160 6276 28172
rect 6328 28160 6334 28212
rect 7006 28160 7012 28212
rect 7064 28200 7070 28212
rect 7653 28203 7711 28209
rect 7653 28200 7665 28203
rect 7064 28172 7665 28200
rect 7064 28160 7070 28172
rect 7653 28169 7665 28172
rect 7699 28169 7711 28203
rect 7653 28163 7711 28169
rect 8386 28160 8392 28212
rect 8444 28160 8450 28212
rect 4816 28132 4844 28160
rect 6104 28132 6132 28160
rect 4448 28104 4844 28132
rect 5934 28104 6132 28132
rect 4448 28076 4476 28104
rect 6546 28092 6552 28144
rect 6604 28132 6610 28144
rect 7101 28135 7159 28141
rect 7101 28132 7113 28135
rect 6604 28104 7113 28132
rect 6604 28092 6610 28104
rect 7101 28101 7113 28104
rect 7147 28101 7159 28135
rect 7101 28095 7159 28101
rect 7193 28135 7251 28141
rect 7193 28101 7205 28135
rect 7239 28132 7251 28135
rect 7239 28104 8248 28132
rect 7239 28101 7251 28104
rect 7193 28095 7251 28101
rect 4430 28024 4436 28076
rect 4488 28024 4494 28076
rect 8220 28073 8248 28104
rect 7837 28067 7895 28073
rect 7837 28064 7849 28067
rect 7576 28036 7849 28064
rect 4706 27956 4712 28008
rect 4764 27956 4770 28008
rect 7009 27999 7067 28005
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 7190 27996 7196 28008
rect 7055 27968 7196 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 7576 27937 7604 28036
rect 7837 28033 7849 28036
rect 7883 28033 7895 28067
rect 7837 28027 7895 28033
rect 8205 28067 8263 28073
rect 8205 28033 8217 28067
rect 8251 28064 8263 28067
rect 8864 28064 8892 28376
rect 8251 28036 8892 28064
rect 8251 28033 8263 28036
rect 8205 28027 8263 28033
rect 7561 27931 7619 27937
rect 7561 27897 7573 27931
rect 7607 27897 7619 27931
rect 7561 27891 7619 27897
rect 1104 27770 8832 27792
rect 1104 27718 2350 27770
rect 2402 27718 2414 27770
rect 2466 27718 2478 27770
rect 2530 27718 2542 27770
rect 2594 27718 2606 27770
rect 2658 27718 7350 27770
rect 7402 27718 7414 27770
rect 7466 27718 7478 27770
rect 7530 27718 7542 27770
rect 7594 27718 7606 27770
rect 7658 27718 8832 27770
rect 1104 27696 8832 27718
rect 8205 27455 8263 27461
rect 8205 27452 8217 27455
rect 7944 27424 8217 27452
rect 7944 27396 7972 27424
rect 8205 27421 8217 27424
rect 8251 27421 8263 27455
rect 8205 27415 8263 27421
rect 8481 27455 8539 27461
rect 8481 27421 8493 27455
rect 8527 27452 8539 27455
rect 8527 27424 8892 27452
rect 8527 27421 8539 27424
rect 8481 27415 8539 27421
rect 7926 27344 7932 27396
rect 7984 27344 7990 27396
rect 8864 27328 8892 27424
rect 7834 27276 7840 27328
rect 7892 27316 7898 27328
rect 8021 27319 8079 27325
rect 8021 27316 8033 27319
rect 7892 27288 8033 27316
rect 7892 27276 7898 27288
rect 8021 27285 8033 27288
rect 8067 27285 8079 27319
rect 8021 27279 8079 27285
rect 8297 27319 8355 27325
rect 8297 27285 8309 27319
rect 8343 27316 8355 27319
rect 8386 27316 8392 27328
rect 8343 27288 8392 27316
rect 8343 27285 8355 27288
rect 8297 27279 8355 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8846 27276 8852 27328
rect 8904 27276 8910 27328
rect 1104 27226 8832 27248
rect 1104 27174 3010 27226
rect 3062 27174 3074 27226
rect 3126 27174 3138 27226
rect 3190 27174 3202 27226
rect 3254 27174 3266 27226
rect 3318 27174 8010 27226
rect 8062 27174 8074 27226
rect 8126 27174 8138 27226
rect 8190 27174 8202 27226
rect 8254 27174 8266 27226
rect 8318 27174 8832 27226
rect 1104 27152 8832 27174
rect 8386 27072 8392 27124
rect 8444 27072 8450 27124
rect 7653 27047 7711 27053
rect 7653 27013 7665 27047
rect 7699 27044 7711 27047
rect 8404 27044 8432 27072
rect 7699 27016 8432 27044
rect 7699 27013 7711 27016
rect 7653 27007 7711 27013
rect 7190 26976 7196 26988
rect 6196 26948 7196 26976
rect 6196 26920 6224 26948
rect 7190 26936 7196 26948
rect 7248 26976 7254 26988
rect 7248 26948 7512 26976
rect 7248 26936 7254 26948
rect 5718 26868 5724 26920
rect 5776 26908 5782 26920
rect 6178 26908 6184 26920
rect 5776 26880 6184 26908
rect 5776 26868 5782 26880
rect 6178 26868 6184 26880
rect 6236 26868 6242 26920
rect 6914 26868 6920 26920
rect 6972 26868 6978 26920
rect 7484 26917 7512 26948
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 8389 26979 8447 26985
rect 8389 26976 8401 26979
rect 8128 26948 8401 26976
rect 7469 26911 7527 26917
rect 7469 26877 7481 26911
rect 7515 26877 7527 26911
rect 7469 26871 7527 26877
rect 8128 26849 8156 26948
rect 8389 26945 8401 26948
rect 8435 26945 8447 26979
rect 8389 26939 8447 26945
rect 8113 26843 8171 26849
rect 8113 26809 8125 26843
rect 8159 26809 8171 26843
rect 8113 26803 8171 26809
rect 6362 26732 6368 26784
rect 6420 26732 6426 26784
rect 7926 26732 7932 26784
rect 7984 26772 7990 26784
rect 8205 26775 8263 26781
rect 8205 26772 8217 26775
rect 7984 26744 8217 26772
rect 7984 26732 7990 26744
rect 8205 26741 8217 26744
rect 8251 26741 8263 26775
rect 8205 26735 8263 26741
rect 1104 26682 8832 26704
rect 1104 26630 2350 26682
rect 2402 26630 2414 26682
rect 2466 26630 2478 26682
rect 2530 26630 2542 26682
rect 2594 26630 2606 26682
rect 2658 26630 7350 26682
rect 7402 26630 7414 26682
rect 7466 26630 7478 26682
rect 7530 26630 7542 26682
rect 7594 26630 7606 26682
rect 7658 26630 8832 26682
rect 1104 26608 8832 26630
rect 4328 26571 4386 26577
rect 4328 26537 4340 26571
rect 4374 26568 4386 26571
rect 5718 26568 5724 26580
rect 4374 26540 5724 26568
rect 4374 26537 4386 26540
rect 4328 26531 4386 26537
rect 5718 26528 5724 26540
rect 5776 26528 5782 26580
rect 5813 26571 5871 26577
rect 5813 26537 5825 26571
rect 5859 26568 5871 26571
rect 6914 26568 6920 26580
rect 5859 26540 6920 26568
rect 5859 26537 5871 26540
rect 5813 26531 5871 26537
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 7742 26528 7748 26580
rect 7800 26528 7806 26580
rect 4065 26435 4123 26441
rect 4065 26401 4077 26435
rect 4111 26432 4123 26435
rect 4430 26432 4436 26444
rect 4111 26404 4436 26432
rect 4111 26401 4123 26404
rect 4065 26395 4123 26401
rect 4430 26392 4436 26404
rect 4488 26392 4494 26444
rect 5905 26435 5963 26441
rect 5905 26401 5917 26435
rect 5951 26432 5963 26435
rect 6730 26432 6736 26444
rect 5951 26404 6736 26432
rect 5951 26401 5963 26404
rect 5905 26395 5963 26401
rect 6730 26392 6736 26404
rect 6788 26392 6794 26444
rect 6914 26392 6920 26444
rect 6972 26432 6978 26444
rect 7653 26435 7711 26441
rect 6972 26404 7328 26432
rect 6972 26392 6978 26404
rect 5566 26268 6132 26296
rect 6104 26228 6132 26268
rect 6178 26256 6184 26308
rect 6236 26256 6242 26308
rect 7300 26228 7328 26404
rect 7653 26401 7665 26435
rect 7699 26432 7711 26435
rect 8297 26435 8355 26441
rect 8297 26432 8309 26435
rect 7699 26404 8309 26432
rect 7699 26401 7711 26404
rect 7653 26395 7711 26401
rect 8297 26401 8309 26404
rect 8343 26401 8355 26435
rect 8297 26395 8355 26401
rect 7742 26324 7748 26376
rect 7800 26364 7806 26376
rect 8018 26364 8024 26376
rect 7800 26336 8024 26364
rect 7800 26324 7806 26336
rect 8018 26324 8024 26336
rect 8076 26324 8082 26376
rect 6104 26200 7328 26228
rect 1104 26138 8832 26160
rect 1104 26086 3010 26138
rect 3062 26086 3074 26138
rect 3126 26086 3138 26138
rect 3190 26086 3202 26138
rect 3254 26086 3266 26138
rect 3318 26086 8010 26138
rect 8062 26086 8074 26138
rect 8126 26086 8138 26138
rect 8190 26086 8202 26138
rect 8254 26086 8266 26138
rect 8318 26086 8832 26138
rect 1104 26064 8832 26086
rect 6086 25984 6092 26036
rect 6144 25984 6150 26036
rect 6178 25984 6184 26036
rect 6236 26024 6242 26036
rect 6365 26027 6423 26033
rect 6365 26024 6377 26027
rect 6236 25996 6377 26024
rect 6236 25984 6242 25996
rect 6365 25993 6377 25996
rect 6411 25993 6423 26027
rect 6365 25987 6423 25993
rect 7926 25984 7932 26036
rect 7984 26024 7990 26036
rect 7984 25996 8156 26024
rect 7984 25984 7990 25996
rect 5721 25959 5779 25965
rect 5721 25925 5733 25959
rect 5767 25956 5779 25959
rect 6104 25956 6132 25984
rect 8128 25965 8156 25996
rect 5767 25928 6132 25956
rect 8113 25959 8171 25965
rect 5767 25925 5779 25928
rect 5721 25919 5779 25925
rect 8113 25925 8125 25959
rect 8159 25925 8171 25959
rect 8113 25919 8171 25925
rect 6549 25891 6607 25897
rect 6549 25888 6561 25891
rect 6196 25860 6561 25888
rect 6196 25829 6224 25860
rect 6549 25857 6561 25860
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 7006 25848 7012 25900
rect 7064 25848 7070 25900
rect 6181 25823 6239 25829
rect 6181 25789 6193 25823
rect 6227 25789 6239 25823
rect 6181 25783 6239 25789
rect 8389 25823 8447 25829
rect 8389 25789 8401 25823
rect 8435 25789 8447 25823
rect 8389 25783 8447 25789
rect 6089 25755 6147 25761
rect 6089 25721 6101 25755
rect 6135 25752 6147 25755
rect 6362 25752 6368 25764
rect 6135 25724 6368 25752
rect 6135 25721 6147 25724
rect 6089 25715 6147 25721
rect 6362 25712 6368 25724
rect 6420 25712 6426 25764
rect 6638 25644 6644 25696
rect 6696 25644 6702 25696
rect 6730 25644 6736 25696
rect 6788 25684 6794 25696
rect 8404 25684 8432 25783
rect 6788 25656 8432 25684
rect 6788 25644 6794 25656
rect 1104 25594 8832 25616
rect 1104 25542 2350 25594
rect 2402 25542 2414 25594
rect 2466 25542 2478 25594
rect 2530 25542 2542 25594
rect 2594 25542 2606 25594
rect 2658 25542 7350 25594
rect 7402 25542 7414 25594
rect 7466 25542 7478 25594
rect 7530 25542 7542 25594
rect 7594 25542 7606 25594
rect 7658 25542 8832 25594
rect 1104 25520 8832 25542
rect 6638 25440 6644 25492
rect 6696 25440 6702 25492
rect 7190 25440 7196 25492
rect 7248 25480 7254 25492
rect 7248 25452 8340 25480
rect 7248 25440 7254 25452
rect 6656 25344 6684 25440
rect 7009 25347 7067 25353
rect 7009 25344 7021 25347
rect 6656 25316 7021 25344
rect 7009 25313 7021 25316
rect 7055 25313 7067 25347
rect 7009 25307 7067 25313
rect 7834 25304 7840 25356
rect 7892 25344 7898 25356
rect 8312 25353 8340 25452
rect 8205 25347 8263 25353
rect 8205 25344 8217 25347
rect 7892 25316 8217 25344
rect 7892 25304 7898 25316
rect 8205 25313 8217 25316
rect 8251 25313 8263 25347
rect 8205 25307 8263 25313
rect 8297 25347 8355 25353
rect 8297 25313 8309 25347
rect 8343 25313 8355 25347
rect 8297 25307 8355 25313
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25245 6975 25279
rect 6917 25239 6975 25245
rect 6638 25100 6644 25152
rect 6696 25140 6702 25152
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 6696 25112 6745 25140
rect 6696 25100 6702 25112
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 6932 25140 6960 25239
rect 7653 25211 7711 25217
rect 7653 25177 7665 25211
rect 7699 25208 7711 25211
rect 8113 25211 8171 25217
rect 8113 25208 8125 25211
rect 7699 25180 8125 25208
rect 7699 25177 7711 25180
rect 7653 25171 7711 25177
rect 8113 25177 8125 25180
rect 8159 25177 8171 25211
rect 8113 25171 8171 25177
rect 7745 25143 7803 25149
rect 7745 25140 7757 25143
rect 6932 25112 7757 25140
rect 6733 25103 6791 25109
rect 7745 25109 7757 25112
rect 7791 25109 7803 25143
rect 7745 25103 7803 25109
rect 1104 25050 8832 25072
rect 1104 24998 3010 25050
rect 3062 24998 3074 25050
rect 3126 24998 3138 25050
rect 3190 24998 3202 25050
rect 3254 24998 3266 25050
rect 3318 24998 8010 25050
rect 8062 24998 8074 25050
rect 8126 24998 8138 25050
rect 8190 24998 8202 25050
rect 8254 24998 8266 25050
rect 8318 24998 8832 25050
rect 1104 24976 8832 24998
rect 6730 24896 6736 24948
rect 6788 24896 6794 24948
rect 7006 24896 7012 24948
rect 7064 24896 7070 24948
rect 6748 24868 6776 24896
rect 6564 24840 6776 24868
rect 7024 24868 7052 24896
rect 7024 24840 7314 24868
rect 6564 24809 6592 24840
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 6656 24704 6837 24732
rect 6656 24608 6684 24704
rect 6825 24701 6837 24704
rect 6871 24701 6883 24735
rect 6825 24695 6883 24701
rect 6638 24556 6644 24608
rect 6696 24556 6702 24608
rect 8297 24599 8355 24605
rect 8297 24565 8309 24599
rect 8343 24596 8355 24599
rect 8386 24596 8392 24608
rect 8343 24568 8392 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 8386 24556 8392 24568
rect 8444 24556 8450 24608
rect 1104 24506 8832 24528
rect 1104 24454 2350 24506
rect 2402 24454 2414 24506
rect 2466 24454 2478 24506
rect 2530 24454 2542 24506
rect 2594 24454 2606 24506
rect 2658 24454 7350 24506
rect 7402 24454 7414 24506
rect 7466 24454 7478 24506
rect 7530 24454 7542 24506
rect 7594 24454 7606 24506
rect 7658 24454 8832 24506
rect 1104 24432 8832 24454
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 7377 24395 7435 24401
rect 7377 24392 7389 24395
rect 7248 24364 7389 24392
rect 7248 24352 7254 24364
rect 7377 24361 7389 24364
rect 7423 24361 7435 24395
rect 7377 24355 7435 24361
rect 7392 24256 7420 24355
rect 8297 24259 8355 24265
rect 8297 24256 8309 24259
rect 7392 24228 8309 24256
rect 8297 24225 8309 24228
rect 8343 24225 8355 24259
rect 8297 24219 8355 24225
rect 5994 24148 6000 24200
rect 6052 24188 6058 24200
rect 6730 24188 6736 24200
rect 6052 24160 6736 24188
rect 6052 24148 6058 24160
rect 6730 24148 6736 24160
rect 6788 24188 6794 24200
rect 7285 24191 7343 24197
rect 7285 24188 7297 24191
rect 6788 24160 7297 24188
rect 6788 24148 6794 24160
rect 7285 24157 7297 24160
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7926 24080 7932 24132
rect 7984 24120 7990 24132
rect 8205 24123 8263 24129
rect 8205 24120 8217 24123
rect 7984 24092 8217 24120
rect 7984 24080 7990 24092
rect 8205 24089 8217 24092
rect 8251 24089 8263 24123
rect 8205 24083 8263 24089
rect 7742 24012 7748 24064
rect 7800 24012 7806 24064
rect 7834 24012 7840 24064
rect 7892 24052 7898 24064
rect 8113 24055 8171 24061
rect 8113 24052 8125 24055
rect 7892 24024 8125 24052
rect 7892 24012 7898 24024
rect 8113 24021 8125 24024
rect 8159 24021 8171 24055
rect 8113 24015 8171 24021
rect 1104 23962 8832 23984
rect 1104 23910 3010 23962
rect 3062 23910 3074 23962
rect 3126 23910 3138 23962
rect 3190 23910 3202 23962
rect 3254 23910 3266 23962
rect 3318 23910 8010 23962
rect 8062 23910 8074 23962
rect 8126 23910 8138 23962
rect 8190 23910 8202 23962
rect 8254 23910 8266 23962
rect 8318 23910 8832 23962
rect 1104 23888 8832 23910
rect 7742 23808 7748 23860
rect 7800 23808 7806 23860
rect 7834 23808 7840 23860
rect 7892 23808 7898 23860
rect 8386 23808 8392 23860
rect 8444 23808 8450 23860
rect 7760 23780 7788 23808
rect 6472 23752 7788 23780
rect 6472 23721 6500 23752
rect 8404 23721 8432 23808
rect 6457 23715 6515 23721
rect 6457 23681 6469 23715
rect 6503 23681 6515 23715
rect 6457 23675 6515 23681
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23681 8447 23715
rect 8389 23675 8447 23681
rect 6840 23644 6868 23675
rect 6472 23616 6868 23644
rect 7193 23647 7251 23653
rect 6472 23588 6500 23616
rect 7193 23613 7205 23647
rect 7239 23644 7251 23647
rect 8294 23644 8300 23656
rect 7239 23616 8300 23644
rect 7239 23613 7251 23616
rect 7193 23607 7251 23613
rect 8294 23604 8300 23616
rect 8352 23604 8358 23656
rect 6454 23536 6460 23588
rect 6512 23536 6518 23588
rect 7009 23579 7067 23585
rect 7009 23545 7021 23579
rect 7055 23576 7067 23579
rect 7098 23576 7104 23588
rect 7055 23548 7104 23576
rect 7055 23545 7067 23548
rect 7009 23539 7067 23545
rect 7098 23536 7104 23548
rect 7156 23536 7162 23588
rect 6641 23511 6699 23517
rect 6641 23477 6653 23511
rect 6687 23508 6699 23511
rect 6730 23508 6736 23520
rect 6687 23480 6736 23508
rect 6687 23477 6699 23480
rect 6641 23471 6699 23477
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 7745 23511 7803 23517
rect 7745 23477 7757 23511
rect 7791 23508 7803 23511
rect 7834 23508 7840 23520
rect 7791 23480 7840 23508
rect 7791 23477 7803 23480
rect 7745 23471 7803 23477
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 1104 23418 8832 23440
rect 1104 23366 2350 23418
rect 2402 23366 2414 23418
rect 2466 23366 2478 23418
rect 2530 23366 2542 23418
rect 2594 23366 2606 23418
rect 2658 23366 7350 23418
rect 7402 23366 7414 23418
rect 7466 23366 7478 23418
rect 7530 23366 7542 23418
rect 7594 23366 7606 23418
rect 7658 23366 8832 23418
rect 1104 23344 8832 23366
rect 8294 23264 8300 23316
rect 8352 23264 8358 23316
rect 6546 23060 6552 23112
rect 6604 23060 6610 23112
rect 6730 22992 6736 23044
rect 6788 23032 6794 23044
rect 6825 23035 6883 23041
rect 6825 23032 6837 23035
rect 6788 23004 6837 23032
rect 6788 22992 6794 23004
rect 6825 23001 6837 23004
rect 6871 23001 6883 23035
rect 6825 22995 6883 23001
rect 6914 22992 6920 23044
rect 6972 23032 6978 23044
rect 7098 23032 7104 23044
rect 6972 23004 7104 23032
rect 6972 22992 6978 23004
rect 7098 22992 7104 23004
rect 7156 23032 7162 23044
rect 7156 23004 7314 23032
rect 7156 22992 7162 23004
rect 1104 22874 8832 22896
rect 1104 22822 3010 22874
rect 3062 22822 3074 22874
rect 3126 22822 3138 22874
rect 3190 22822 3202 22874
rect 3254 22822 3266 22874
rect 3318 22822 8010 22874
rect 8062 22822 8074 22874
rect 8126 22822 8138 22874
rect 8190 22822 8202 22874
rect 8254 22822 8266 22874
rect 8318 22822 8832 22874
rect 1104 22800 8832 22822
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 7208 22732 7757 22760
rect 7208 22633 7236 22732
rect 7745 22729 7757 22732
rect 7791 22729 7803 22763
rect 7745 22723 7803 22729
rect 7834 22720 7840 22772
rect 7892 22760 7898 22772
rect 8113 22763 8171 22769
rect 8113 22760 8125 22763
rect 7892 22732 8125 22760
rect 7892 22720 7898 22732
rect 8113 22729 8125 22732
rect 8159 22729 8171 22763
rect 8113 22723 8171 22729
rect 8386 22720 8392 22772
rect 8444 22720 8450 22772
rect 7374 22652 7380 22704
rect 7432 22692 7438 22704
rect 8205 22695 8263 22701
rect 8205 22692 8217 22695
rect 7432 22664 8217 22692
rect 7432 22652 7438 22664
rect 8205 22661 8217 22664
rect 8251 22661 8263 22695
rect 8205 22655 8263 22661
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 6932 22556 6960 22587
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 7340 22596 7481 22624
rect 7340 22584 7346 22596
rect 7469 22593 7481 22596
rect 7515 22593 7527 22627
rect 8404 22624 8432 22720
rect 7469 22587 7527 22593
rect 7576 22596 8432 22624
rect 7576 22556 7604 22596
rect 6932 22528 7604 22556
rect 8297 22559 8355 22565
rect 8297 22525 8309 22559
rect 8343 22525 8355 22559
rect 8297 22519 8355 22525
rect 7653 22491 7711 22497
rect 7653 22457 7665 22491
rect 7699 22488 7711 22491
rect 7834 22488 7840 22500
rect 7699 22460 7840 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 7834 22448 7840 22460
rect 7892 22448 7898 22500
rect 7926 22448 7932 22500
rect 7984 22488 7990 22500
rect 8312 22488 8340 22519
rect 7984 22460 8340 22488
rect 7984 22448 7990 22460
rect 6638 22380 6644 22432
rect 6696 22420 6702 22432
rect 7006 22420 7012 22432
rect 6696 22392 7012 22420
rect 6696 22380 6702 22392
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 7101 22423 7159 22429
rect 7101 22389 7113 22423
rect 7147 22420 7159 22423
rect 7282 22420 7288 22432
rect 7147 22392 7288 22420
rect 7147 22389 7159 22392
rect 7101 22383 7159 22389
rect 7282 22380 7288 22392
rect 7340 22380 7346 22432
rect 7377 22423 7435 22429
rect 7377 22389 7389 22423
rect 7423 22420 7435 22423
rect 7742 22420 7748 22432
rect 7423 22392 7748 22420
rect 7423 22389 7435 22392
rect 7377 22383 7435 22389
rect 7742 22380 7748 22392
rect 7800 22380 7806 22432
rect 1104 22330 8832 22352
rect 1104 22278 2350 22330
rect 2402 22278 2414 22330
rect 2466 22278 2478 22330
rect 2530 22278 2542 22330
rect 2594 22278 2606 22330
rect 2658 22278 7350 22330
rect 7402 22278 7414 22330
rect 7466 22278 7478 22330
rect 7530 22278 7542 22330
rect 7594 22278 7606 22330
rect 7658 22278 8832 22330
rect 1104 22256 8832 22278
rect 6546 22040 6552 22092
rect 6604 22080 6610 22092
rect 8297 22083 8355 22089
rect 8297 22080 8309 22083
rect 6604 22052 8309 22080
rect 6604 22040 6610 22052
rect 8297 22049 8309 22052
rect 8343 22049 8355 22083
rect 8297 22043 8355 22049
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 7742 21904 7748 21956
rect 7800 21944 7806 21956
rect 8021 21947 8079 21953
rect 8021 21944 8033 21947
rect 7800 21916 8033 21944
rect 7800 21904 7806 21916
rect 8021 21913 8033 21916
rect 8067 21913 8079 21947
rect 8021 21907 8079 21913
rect 6549 21879 6607 21885
rect 6549 21845 6561 21879
rect 6595 21876 6607 21879
rect 7006 21876 7012 21888
rect 6595 21848 7012 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 7006 21836 7012 21848
rect 7064 21836 7070 21888
rect 1104 21786 8832 21808
rect 1104 21734 3010 21786
rect 3062 21734 3074 21786
rect 3126 21734 3138 21786
rect 3190 21734 3202 21786
rect 3254 21734 3266 21786
rect 3318 21734 8010 21786
rect 8062 21734 8074 21786
rect 8126 21734 8138 21786
rect 8190 21734 8202 21786
rect 8254 21734 8266 21786
rect 8318 21734 8832 21786
rect 1104 21712 8832 21734
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 8205 21675 8263 21681
rect 8205 21672 8217 21675
rect 6963 21644 8217 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 8205 21641 8217 21644
rect 8251 21641 8263 21675
rect 8205 21635 8263 21641
rect 8294 21604 8300 21616
rect 6748 21576 8300 21604
rect 6748 21545 6776 21576
rect 8294 21564 8300 21576
rect 8352 21564 8358 21616
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 7006 21496 7012 21548
rect 7064 21496 7070 21548
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21536 7711 21539
rect 8113 21539 8171 21545
rect 8113 21536 8125 21539
rect 7699 21508 8125 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 8113 21505 8125 21508
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 7926 21428 7932 21480
rect 7984 21468 7990 21480
rect 8297 21471 8355 21477
rect 8297 21468 8309 21471
rect 7984 21440 8309 21468
rect 7984 21428 7990 21440
rect 8297 21437 8309 21440
rect 8343 21437 8355 21471
rect 8297 21431 8355 21437
rect 7742 21292 7748 21344
rect 7800 21292 7806 21344
rect 1104 21242 8832 21264
rect 1104 21190 2350 21242
rect 2402 21190 2414 21242
rect 2466 21190 2478 21242
rect 2530 21190 2542 21242
rect 2594 21190 2606 21242
rect 2658 21190 7350 21242
rect 7402 21190 7414 21242
rect 7466 21190 7478 21242
rect 7530 21190 7542 21242
rect 7594 21190 7606 21242
rect 7658 21190 8832 21242
rect 1104 21168 8832 21190
rect 6914 21088 6920 21140
rect 6972 21128 6978 21140
rect 7282 21128 7288 21140
rect 6972 21100 7288 21128
rect 6972 21088 6978 21100
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 6546 20952 6552 21004
rect 6604 20952 6610 21004
rect 6825 20859 6883 20865
rect 6825 20825 6837 20859
rect 6871 20856 6883 20859
rect 7098 20856 7104 20868
rect 6871 20828 7104 20856
rect 6871 20825 6883 20828
rect 6825 20819 6883 20825
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 7282 20816 7288 20868
rect 7340 20816 7346 20868
rect 8297 20791 8355 20797
rect 8297 20757 8309 20791
rect 8343 20788 8355 20791
rect 8386 20788 8392 20800
rect 8343 20760 8392 20788
rect 8343 20757 8355 20760
rect 8297 20751 8355 20757
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 1104 20698 8832 20720
rect 1104 20646 3010 20698
rect 3062 20646 3074 20698
rect 3126 20646 3138 20698
rect 3190 20646 3202 20698
rect 3254 20646 3266 20698
rect 3318 20646 8010 20698
rect 8062 20646 8074 20698
rect 8126 20646 8138 20698
rect 8190 20646 8202 20698
rect 8254 20646 8266 20698
rect 8318 20646 8832 20698
rect 1104 20624 8832 20646
rect 7098 20544 7104 20596
rect 7156 20584 7162 20596
rect 7193 20587 7251 20593
rect 7193 20584 7205 20587
rect 7156 20556 7205 20584
rect 7156 20544 7162 20556
rect 7193 20553 7205 20556
rect 7239 20553 7251 20587
rect 7193 20547 7251 20553
rect 7742 20544 7748 20596
rect 7800 20544 7806 20596
rect 7926 20544 7932 20596
rect 7984 20584 7990 20596
rect 7984 20556 8248 20584
rect 7984 20544 7990 20556
rect 7760 20516 7788 20544
rect 8220 20528 8248 20556
rect 7392 20488 7788 20516
rect 7392 20457 7420 20488
rect 8202 20476 8208 20528
rect 8260 20476 8266 20528
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20448 7527 20451
rect 7926 20448 7932 20460
rect 7515 20420 7932 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 8110 20408 8116 20460
rect 8168 20408 8174 20460
rect 8220 20448 8248 20476
rect 8220 20420 8340 20448
rect 7190 20340 7196 20392
rect 7248 20380 7254 20392
rect 8312 20389 8340 20420
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 7248 20352 8217 20380
rect 7248 20340 7254 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 8205 20343 8263 20349
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 7653 20315 7711 20321
rect 7653 20281 7665 20315
rect 7699 20312 7711 20315
rect 7834 20312 7840 20324
rect 7699 20284 7840 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 7834 20272 7840 20284
rect 7892 20272 7898 20324
rect 7098 20204 7104 20256
rect 7156 20244 7162 20256
rect 7282 20244 7288 20256
rect 7156 20216 7288 20244
rect 7156 20204 7162 20216
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7742 20204 7748 20256
rect 7800 20204 7806 20256
rect 1104 20154 8832 20176
rect 1104 20102 2350 20154
rect 2402 20102 2414 20154
rect 2466 20102 2478 20154
rect 2530 20102 2542 20154
rect 2594 20102 2606 20154
rect 2658 20102 7350 20154
rect 7402 20102 7414 20154
rect 7466 20102 7478 20154
rect 7530 20102 7542 20154
rect 7594 20102 7606 20154
rect 7658 20102 8832 20154
rect 1104 20080 8832 20102
rect 7742 20000 7748 20052
rect 7800 20000 7806 20052
rect 7837 20043 7895 20049
rect 7837 20009 7849 20043
rect 7883 20040 7895 20043
rect 8110 20040 8116 20052
rect 7883 20012 8116 20040
rect 7883 20009 7895 20012
rect 7837 20003 7895 20009
rect 8110 20000 8116 20012
rect 8168 20000 8174 20052
rect 6730 19932 6736 19984
rect 6788 19972 6794 19984
rect 6825 19975 6883 19981
rect 6825 19972 6837 19975
rect 6788 19944 6837 19972
rect 6788 19932 6794 19944
rect 6825 19941 6837 19944
rect 6871 19941 6883 19975
rect 6825 19935 6883 19941
rect 7760 19904 7788 20000
rect 7024 19876 7788 19904
rect 7024 19845 7052 19876
rect 8386 19864 8392 19916
rect 8444 19864 8450 19916
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19836 7251 19839
rect 7239 19808 8892 19836
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 6564 19768 6592 19799
rect 8294 19768 8300 19780
rect 6564 19740 8300 19768
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 6733 19703 6791 19709
rect 6733 19669 6745 19703
rect 6779 19700 6791 19703
rect 7190 19700 7196 19712
rect 6779 19672 7196 19700
rect 6779 19669 6791 19672
rect 6733 19663 6791 19669
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 7745 19703 7803 19709
rect 7745 19669 7757 19703
rect 7791 19700 7803 19703
rect 7834 19700 7840 19712
rect 7791 19672 7840 19700
rect 7791 19669 7803 19672
rect 7745 19663 7803 19669
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 8202 19660 8208 19712
rect 8260 19700 8266 19712
rect 8386 19700 8392 19712
rect 8260 19672 8392 19700
rect 8260 19660 8266 19672
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 1104 19610 8832 19632
rect 1104 19558 3010 19610
rect 3062 19558 3074 19610
rect 3126 19558 3138 19610
rect 3190 19558 3202 19610
rect 3254 19558 3266 19610
rect 3318 19558 8010 19610
rect 8062 19558 8074 19610
rect 8126 19558 8138 19610
rect 8190 19558 8202 19610
rect 8254 19558 8266 19610
rect 8318 19558 8832 19610
rect 1104 19536 8832 19558
rect 7190 19456 7196 19508
rect 7248 19456 7254 19508
rect 8297 19499 8355 19505
rect 8297 19465 8309 19499
rect 8343 19496 8355 19499
rect 8864 19496 8892 19808
rect 8343 19468 8892 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 6730 19388 6736 19440
rect 6788 19428 6794 19440
rect 6825 19431 6883 19437
rect 6825 19428 6837 19431
rect 6788 19400 6837 19428
rect 6788 19388 6794 19400
rect 6825 19397 6837 19400
rect 6871 19397 6883 19431
rect 7208 19428 7236 19456
rect 7208 19400 7314 19428
rect 6825 19391 6883 19397
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 1104 19066 8832 19088
rect 1104 19014 2350 19066
rect 2402 19014 2414 19066
rect 2466 19014 2478 19066
rect 2530 19014 2542 19066
rect 2594 19014 2606 19066
rect 2658 19014 7350 19066
rect 7402 19014 7414 19066
rect 7466 19014 7478 19066
rect 7530 19014 7542 19066
rect 7594 19014 7606 19066
rect 7658 19014 8832 19066
rect 1104 18992 8832 19014
rect 8202 18912 8208 18964
rect 8260 18912 8266 18964
rect 7926 18844 7932 18896
rect 7984 18884 7990 18896
rect 8220 18884 8248 18912
rect 7984 18856 8340 18884
rect 7984 18844 7990 18856
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 8312 18825 8340 18856
rect 8205 18819 8263 18825
rect 8205 18816 8217 18819
rect 7800 18788 8217 18816
rect 7800 18776 7806 18788
rect 8205 18785 8217 18788
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 8297 18819 8355 18825
rect 8297 18785 8309 18819
rect 8343 18785 8355 18819
rect 8297 18779 8355 18785
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18748 7435 18751
rect 7423 18720 7788 18748
rect 7423 18717 7435 18720
rect 7377 18711 7435 18717
rect 7190 18572 7196 18624
rect 7248 18572 7254 18624
rect 7760 18621 7788 18720
rect 7834 18708 7840 18760
rect 7892 18748 7898 18760
rect 8113 18751 8171 18757
rect 8113 18748 8125 18751
rect 7892 18720 8125 18748
rect 7892 18708 7898 18720
rect 8113 18717 8125 18720
rect 8159 18717 8171 18751
rect 8113 18711 8171 18717
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18581 7803 18615
rect 7745 18575 7803 18581
rect 1104 18522 8832 18544
rect 1104 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 3202 18522
rect 3254 18470 3266 18522
rect 3318 18470 8010 18522
rect 8062 18470 8074 18522
rect 8126 18470 8138 18522
rect 8190 18470 8202 18522
rect 8254 18470 8266 18522
rect 8318 18470 8832 18522
rect 1104 18448 8832 18470
rect 7190 18408 7196 18420
rect 6840 18380 7196 18408
rect 6840 18349 6868 18380
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18309 6883 18343
rect 6825 18303 6883 18309
rect 6546 18232 6552 18284
rect 6604 18232 6610 18284
rect 7926 18232 7932 18284
rect 7984 18232 7990 18284
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7944 18204 7972 18232
rect 7340 18176 7972 18204
rect 7340 18164 7346 18176
rect 8297 18071 8355 18077
rect 8297 18037 8309 18071
rect 8343 18068 8355 18071
rect 8386 18068 8392 18080
rect 8343 18040 8392 18068
rect 8343 18037 8355 18040
rect 8297 18031 8355 18037
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 1104 17978 8832 18000
rect 1104 17926 2350 17978
rect 2402 17926 2414 17978
rect 2466 17926 2478 17978
rect 2530 17926 2542 17978
rect 2594 17926 2606 17978
rect 2658 17926 7350 17978
rect 7402 17926 7414 17978
rect 7466 17926 7478 17978
rect 7530 17926 7542 17978
rect 7594 17926 7606 17978
rect 7658 17926 8832 17978
rect 1104 17904 8832 17926
rect 7834 17864 7840 17876
rect 7668 17836 7840 17864
rect 7668 17805 7696 17836
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 7285 17799 7343 17805
rect 7285 17765 7297 17799
rect 7331 17765 7343 17799
rect 7285 17759 7343 17765
rect 7653 17799 7711 17805
rect 7653 17765 7665 17799
rect 7699 17796 7711 17799
rect 7699 17768 8340 17796
rect 7699 17765 7711 17768
rect 7653 17759 7711 17765
rect 7300 17728 7328 17759
rect 8312 17737 8340 17768
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 7300 17700 8217 17728
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 7147 17632 8524 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 8496 17604 8524 17632
rect 6914 17552 6920 17604
rect 6972 17592 6978 17604
rect 7469 17595 7527 17601
rect 7469 17592 7481 17595
rect 6972 17564 7481 17592
rect 6972 17552 6978 17564
rect 7116 17536 7144 17564
rect 7469 17561 7481 17564
rect 7515 17561 7527 17595
rect 7469 17555 7527 17561
rect 8478 17552 8484 17604
rect 8536 17552 8542 17604
rect 7098 17484 7104 17536
rect 7156 17484 7162 17536
rect 7742 17484 7748 17536
rect 7800 17484 7806 17536
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7892 17496 8125 17524
rect 7892 17484 7898 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 1104 17434 8832 17456
rect 1104 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 3202 17434
rect 3254 17382 3266 17434
rect 3318 17382 8010 17434
rect 8062 17382 8074 17434
rect 8126 17382 8138 17434
rect 8190 17382 8202 17434
rect 8254 17382 8266 17434
rect 8318 17382 8832 17434
rect 1104 17360 8832 17382
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 7834 17280 7840 17332
rect 7892 17280 7898 17332
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 7009 17187 7067 17193
rect 6595 17156 6776 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6748 17128 6776 17156
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7760 17184 7788 17280
rect 7055 17156 7788 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 6730 17076 6736 17128
rect 6788 17076 6794 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 8294 17116 8300 17128
rect 7239 17088 8300 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 6696 17020 6837 17048
rect 6696 17008 6702 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 6733 16983 6791 16989
rect 6733 16949 6745 16983
rect 6779 16980 6791 16983
rect 6914 16980 6920 16992
rect 6779 16952 6920 16980
rect 6779 16949 6791 16952
rect 6733 16943 6791 16949
rect 6914 16940 6920 16952
rect 6972 16940 6978 16992
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16980 7803 16983
rect 7926 16980 7932 16992
rect 7791 16952 7932 16980
rect 7791 16949 7803 16952
rect 7745 16943 7803 16949
rect 7926 16940 7932 16952
rect 7984 16940 7990 16992
rect 1104 16890 8832 16912
rect 1104 16838 2350 16890
rect 2402 16838 2414 16890
rect 2466 16838 2478 16890
rect 2530 16838 2542 16890
rect 2594 16838 2606 16890
rect 2658 16838 7350 16890
rect 7402 16838 7414 16890
rect 7466 16838 7478 16890
rect 7530 16838 7542 16890
rect 7594 16838 7606 16890
rect 7658 16838 8832 16890
rect 1104 16816 8832 16838
rect 6638 16736 6644 16788
rect 6696 16736 6702 16788
rect 8294 16736 8300 16788
rect 8352 16736 8358 16788
rect 6546 16600 6552 16652
rect 6604 16600 6610 16652
rect 6656 16640 6684 16736
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6656 16612 6837 16640
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 7834 16464 7840 16516
rect 7892 16464 7898 16516
rect 1104 16346 8832 16368
rect 1104 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 3202 16346
rect 3254 16294 3266 16346
rect 3318 16294 8010 16346
rect 8062 16294 8074 16346
rect 8126 16294 8138 16346
rect 8190 16294 8202 16346
rect 8254 16294 8266 16346
rect 8318 16294 8832 16346
rect 1104 16272 8832 16294
rect 7745 16235 7803 16241
rect 7745 16201 7757 16235
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 6914 16056 6920 16108
rect 6972 16056 6978 16108
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16096 7251 16099
rect 7760 16096 7788 16195
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 8113 16235 8171 16241
rect 8113 16232 8125 16235
rect 7984 16204 8125 16232
rect 7984 16192 7990 16204
rect 8113 16201 8125 16204
rect 8159 16201 8171 16235
rect 8113 16195 8171 16201
rect 7239 16068 7788 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 6932 16028 6960 16056
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 6932 16000 8217 16028
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 7834 15920 7840 15972
rect 7892 15960 7898 15972
rect 8312 15960 8340 15991
rect 7892 15932 8340 15960
rect 7892 15920 7898 15932
rect 7377 15895 7435 15901
rect 7377 15861 7389 15895
rect 7423 15892 7435 15895
rect 7926 15892 7932 15904
rect 7423 15864 7932 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 1104 15802 8832 15824
rect 1104 15750 2350 15802
rect 2402 15750 2414 15802
rect 2466 15750 2478 15802
rect 2530 15750 2542 15802
rect 2594 15750 2606 15802
rect 2658 15750 7350 15802
rect 7402 15750 7414 15802
rect 7466 15750 7478 15802
rect 7530 15750 7542 15802
rect 7594 15750 7606 15802
rect 7658 15750 8832 15802
rect 1104 15728 8832 15750
rect 7926 15512 7932 15564
rect 7984 15552 7990 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7984 15524 8033 15552
rect 7984 15512 7990 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 6914 15444 6920 15496
rect 6972 15444 6978 15496
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8386 15484 8392 15496
rect 8343 15456 8392 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 6638 15348 6644 15360
rect 6595 15320 6644 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 1104 15258 8832 15280
rect 1104 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 3202 15258
rect 3254 15206 3266 15258
rect 3318 15206 8010 15258
rect 8062 15206 8074 15258
rect 8126 15206 8138 15258
rect 8190 15206 8202 15258
rect 8254 15206 8266 15258
rect 8318 15206 8832 15258
rect 1104 15184 8832 15206
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 8386 15144 8392 15156
rect 6604 15116 8392 15144
rect 6604 15104 6610 15116
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 8036 15085 8064 15116
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 7285 15079 7343 15085
rect 7285 15076 7297 15079
rect 6880 15048 7297 15076
rect 6880 15036 6886 15048
rect 7285 15045 7297 15048
rect 7331 15045 7343 15079
rect 7285 15039 7343 15045
rect 8021 15079 8079 15085
rect 8021 15045 8033 15079
rect 8067 15045 8079 15079
rect 8021 15039 8079 15045
rect 6638 14968 6644 15020
rect 6696 14968 6702 15020
rect 8481 15011 8539 15017
rect 8481 14977 8493 15011
rect 8527 15008 8539 15011
rect 8527 14980 8892 15008
rect 8527 14977 8539 14980
rect 8481 14971 8539 14977
rect 8864 14884 8892 14980
rect 8846 14832 8852 14884
rect 8904 14832 8910 14884
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 8260 14776 8309 14804
rect 8260 14764 8266 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8297 14767 8355 14773
rect 1104 14714 8832 14736
rect 1104 14662 2350 14714
rect 2402 14662 2414 14714
rect 2466 14662 2478 14714
rect 2530 14662 2542 14714
rect 2594 14662 2606 14714
rect 2658 14662 7350 14714
rect 7402 14662 7414 14714
rect 7466 14662 7478 14714
rect 7530 14662 7542 14714
rect 7594 14662 7606 14714
rect 7658 14662 8832 14714
rect 1104 14640 8832 14662
rect 6914 14560 6920 14612
rect 6972 14560 6978 14612
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7248 14572 8156 14600
rect 7248 14560 7254 14572
rect 6932 14532 6960 14560
rect 7282 14532 7288 14544
rect 6932 14504 7288 14532
rect 7282 14492 7288 14504
rect 7340 14492 7346 14544
rect 6822 14356 6828 14408
rect 6880 14356 6886 14408
rect 8128 14405 8156 14572
rect 8202 14424 8208 14476
rect 8260 14424 8266 14476
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14396 7159 14399
rect 8113 14399 8171 14405
rect 7147 14368 7788 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 6086 14288 6092 14340
rect 6144 14288 6150 14340
rect 6454 14288 6460 14340
rect 6512 14328 6518 14340
rect 7561 14331 7619 14337
rect 7561 14328 7573 14331
rect 6512 14300 7573 14328
rect 6512 14288 6518 14300
rect 7561 14297 7573 14300
rect 7607 14297 7619 14331
rect 7561 14291 7619 14297
rect 6914 14220 6920 14272
rect 6972 14220 6978 14272
rect 7760 14269 7788 14368
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8312 14396 8340 14427
rect 8113 14359 8171 14365
rect 8220 14368 8340 14396
rect 7745 14263 7803 14269
rect 7745 14229 7757 14263
rect 7791 14229 7803 14263
rect 7745 14223 7803 14229
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8220 14260 8248 14368
rect 7892 14232 8248 14260
rect 7892 14220 7898 14232
rect 1104 14170 8832 14192
rect 1104 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 3202 14170
rect 3254 14118 3266 14170
rect 3318 14118 8010 14170
rect 8062 14118 8074 14170
rect 8126 14118 8138 14170
rect 8190 14118 8202 14170
rect 8254 14118 8266 14170
rect 8318 14118 8832 14170
rect 1104 14096 8832 14118
rect 6825 13991 6883 13997
rect 6825 13957 6837 13991
rect 6871 13988 6883 13991
rect 6914 13988 6920 14000
rect 6871 13960 6920 13988
rect 6871 13957 6883 13960
rect 6825 13951 6883 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7282 13948 7288 14000
rect 7340 13948 7346 14000
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 7892 13824 8309 13852
rect 7892 13812 7898 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 1104 13626 8832 13648
rect 1104 13574 2350 13626
rect 2402 13574 2414 13626
rect 2466 13574 2478 13626
rect 2530 13574 2542 13626
rect 2594 13574 2606 13626
rect 2658 13574 7350 13626
rect 7402 13574 7414 13626
rect 7466 13574 7478 13626
rect 7530 13574 7542 13626
rect 7594 13574 7606 13626
rect 7658 13574 8832 13626
rect 1104 13552 8832 13574
rect 6641 13515 6699 13521
rect 6641 13481 6653 13515
rect 6687 13512 6699 13515
rect 6687 13484 8248 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 7745 13447 7803 13453
rect 7745 13444 7757 13447
rect 6932 13416 7757 13444
rect 6932 13317 6960 13416
rect 7745 13413 7757 13416
rect 7791 13413 7803 13447
rect 7745 13407 7803 13413
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7834 13376 7840 13388
rect 7147 13348 7840 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8220 13385 8248 13484
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13345 8263 13379
rect 8205 13339 8263 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7024 13280 8340 13308
rect 6472 13240 6500 13271
rect 7024 13240 7052 13280
rect 8312 13252 8340 13280
rect 6472 13212 7052 13240
rect 7653 13243 7711 13249
rect 7653 13209 7665 13243
rect 7699 13240 7711 13243
rect 8113 13243 8171 13249
rect 8113 13240 8125 13243
rect 7699 13212 8125 13240
rect 7699 13209 7711 13212
rect 7653 13203 7711 13209
rect 8113 13209 8125 13212
rect 8159 13209 8171 13243
rect 8113 13203 8171 13209
rect 8294 13200 8300 13252
rect 8352 13200 8358 13252
rect 6730 13132 6736 13184
rect 6788 13132 6794 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8404 13172 8432 13339
rect 7892 13144 8432 13172
rect 7892 13132 7898 13144
rect 1104 13082 8832 13104
rect 1104 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 3202 13082
rect 3254 13030 3266 13082
rect 3318 13030 8010 13082
rect 8062 13030 8074 13082
rect 8126 13030 8138 13082
rect 8190 13030 8202 13082
rect 8254 13030 8266 13082
rect 8318 13030 8832 13082
rect 1104 13008 8832 13030
rect 6730 12928 6736 12980
rect 6788 12928 6794 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7190 12968 7196 12980
rect 7064 12940 7196 12968
rect 7064 12928 7070 12940
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 6748 12900 6776 12928
rect 6825 12903 6883 12909
rect 6825 12900 6837 12903
rect 6748 12872 6837 12900
rect 6825 12869 6837 12872
rect 6871 12869 6883 12903
rect 7208 12900 7236 12928
rect 7208 12872 7314 12900
rect 6825 12863 6883 12869
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6546 12832 6552 12844
rect 6144 12804 6552 12832
rect 6144 12792 6150 12804
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 8294 12588 8300 12640
rect 8352 12588 8358 12640
rect 1104 12538 8832 12560
rect 1104 12486 2350 12538
rect 2402 12486 2414 12538
rect 2466 12486 2478 12538
rect 2530 12486 2542 12538
rect 2594 12486 2606 12538
rect 2658 12486 7350 12538
rect 7402 12486 7414 12538
rect 7466 12486 7478 12538
rect 7530 12486 7542 12538
rect 7594 12486 7606 12538
rect 7658 12486 8832 12538
rect 1104 12464 8832 12486
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7892 12260 8309 12288
rect 7892 12248 7898 12260
rect 8297 12257 8309 12260
rect 8343 12288 8355 12291
rect 8570 12288 8576 12300
rect 8343 12260 8576 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 7926 12220 7932 12232
rect 7515 12192 7932 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 6788 12124 8217 12152
rect 6788 12112 6794 12124
rect 8205 12121 8217 12124
rect 8251 12121 8263 12155
rect 8205 12115 8263 12121
rect 7650 12044 7656 12096
rect 7708 12044 7714 12096
rect 7742 12044 7748 12096
rect 7800 12044 7806 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 7892 12056 8125 12084
rect 7892 12044 7898 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 1104 11994 8832 12016
rect 1104 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 3202 11994
rect 3254 11942 3266 11994
rect 3318 11942 8010 11994
rect 8062 11942 8074 11994
rect 8126 11942 8138 11994
rect 8190 11942 8202 11994
rect 8254 11942 8266 11994
rect 8318 11942 8832 11994
rect 1104 11920 8832 11942
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 7742 11840 7748 11892
rect 7800 11840 7806 11892
rect 7834 11840 7840 11892
rect 7892 11840 7898 11892
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7760 11744 7788 11840
rect 7055 11716 7788 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 6564 11608 6592 11707
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 7190 11636 7196 11688
rect 7248 11636 7254 11688
rect 8478 11636 8484 11688
rect 8536 11636 8542 11688
rect 8496 11608 8524 11636
rect 6564 11580 8524 11608
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 7745 11543 7803 11549
rect 7745 11509 7757 11543
rect 7791 11540 7803 11543
rect 7926 11540 7932 11552
rect 7791 11512 7932 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 1104 11450 8832 11472
rect 1104 11398 2350 11450
rect 2402 11398 2414 11450
rect 2466 11398 2478 11450
rect 2530 11398 2542 11450
rect 2594 11398 2606 11450
rect 2658 11398 7350 11450
rect 7402 11398 7414 11450
rect 7466 11398 7478 11450
rect 7530 11398 7542 11450
rect 7594 11398 7606 11450
rect 7658 11398 8832 11450
rect 1104 11376 8832 11398
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 8297 11339 8355 11345
rect 8297 11336 8309 11339
rect 7248 11308 8309 11336
rect 7248 11296 7254 11308
rect 8297 11305 8309 11308
rect 8343 11305 8355 11339
rect 8297 11299 8355 11305
rect 6546 11160 6552 11212
rect 6604 11160 6610 11212
rect 6822 11160 6828 11212
rect 6880 11160 6886 11212
rect 7024 11036 7314 11064
rect 7024 11008 7052 11036
rect 7006 10956 7012 11008
rect 7064 10956 7070 11008
rect 1104 10906 8832 10928
rect 1104 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 3202 10906
rect 3254 10854 3266 10906
rect 3318 10854 8010 10906
rect 8062 10854 8074 10906
rect 8126 10854 8138 10906
rect 8190 10854 8202 10906
rect 8254 10854 8266 10906
rect 8318 10854 8832 10906
rect 1104 10832 8832 10854
rect 7745 10795 7803 10801
rect 7745 10761 7757 10795
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 7760 10656 7788 10755
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7984 10764 8125 10792
rect 7984 10752 7990 10764
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8113 10755 8171 10761
rect 7423 10628 7788 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7800 10560 8217 10588
rect 7800 10548 7806 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8570 10588 8576 10600
rect 8435 10560 8576 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 7190 10412 7196 10464
rect 7248 10412 7254 10464
rect 1104 10362 8832 10384
rect 1104 10310 2350 10362
rect 2402 10310 2414 10362
rect 2466 10310 2478 10362
rect 2530 10310 2542 10362
rect 2594 10310 2606 10362
rect 2658 10310 7350 10362
rect 7402 10310 7414 10362
rect 7466 10310 7478 10362
rect 7530 10310 7542 10362
rect 7594 10310 7606 10362
rect 7658 10310 8832 10362
rect 1104 10288 8832 10310
rect 6546 10072 6552 10124
rect 6604 10072 6610 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7190 10112 7196 10124
rect 6871 10084 7196 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7282 9976 7288 9988
rect 7024 9948 7288 9976
rect 7024 9920 7052 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 7006 9868 7012 9920
rect 7064 9868 7070 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8386 9908 8392 9920
rect 8343 9880 8392 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 1104 9818 8832 9840
rect 1104 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 3202 9818
rect 3254 9766 3266 9818
rect 3318 9766 8010 9818
rect 8062 9766 8074 9818
rect 8126 9766 8138 9818
rect 8190 9766 8202 9818
rect 8254 9766 8266 9818
rect 8318 9766 8832 9818
rect 1104 9744 8832 9766
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7064 9540 7481 9568
rect 7064 9528 7070 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 6788 9472 8217 9500
rect 6788 9460 6794 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8570 9500 8576 9512
rect 8435 9472 8576 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 7653 9435 7711 9441
rect 7653 9401 7665 9435
rect 7699 9432 7711 9435
rect 7834 9432 7840 9444
rect 7699 9404 7840 9432
rect 7699 9401 7711 9404
rect 7653 9395 7711 9401
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 7926 9392 7932 9444
rect 7984 9432 7990 9444
rect 8404 9432 8432 9463
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 7984 9404 8432 9432
rect 7984 9392 7990 9404
rect 7742 9324 7748 9376
rect 7800 9324 7806 9376
rect 1104 9274 8832 9296
rect 1104 9222 2350 9274
rect 2402 9222 2414 9274
rect 2466 9222 2478 9274
rect 2530 9222 2542 9274
rect 2594 9222 2606 9274
rect 2658 9222 7350 9274
rect 7402 9222 7414 9274
rect 7466 9222 7478 9274
rect 7530 9222 7542 9274
rect 7594 9222 7606 9274
rect 7658 9222 8832 9274
rect 1104 9200 8832 9222
rect 6730 9120 6736 9172
rect 6788 9120 6794 9172
rect 7742 9120 7748 9172
rect 7800 9120 7806 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 8110 9160 8116 9172
rect 7883 9132 8116 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 7760 9024 7788 9120
rect 7024 8996 7788 9024
rect 7024 8965 7052 8996
rect 8386 8984 8392 9036
rect 8444 8984 8450 9036
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 6564 8888 6592 8919
rect 7190 8916 7196 8968
rect 7248 8916 7254 8968
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 8312 8888 8340 8916
rect 6564 8860 8340 8888
rect 6822 8780 6828 8832
rect 6880 8780 6886 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 1104 8730 8832 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 8010 8730
rect 8062 8678 8074 8730
rect 8126 8678 8138 8730
rect 8190 8678 8202 8730
rect 8254 8678 8266 8730
rect 8318 8678 8832 8730
rect 1104 8656 8832 8678
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 7248 8588 8309 8616
rect 7248 8576 7254 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 7282 8508 7288 8560
rect 7340 8508 7346 8560
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 5994 8372 6000 8424
rect 6052 8372 6058 8424
rect 6822 8372 6828 8424
rect 6880 8372 6886 8424
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5132 8248 5457 8276
rect 5132 8236 5138 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5445 8239 5503 8245
rect 1104 8186 8832 8208
rect 1104 8134 2350 8186
rect 2402 8134 2414 8186
rect 2466 8134 2478 8186
rect 2530 8134 2542 8186
rect 2594 8134 2606 8186
rect 2658 8134 7350 8186
rect 7402 8134 7414 8186
rect 7466 8134 7478 8186
rect 7530 8134 7542 8186
rect 7594 8134 7606 8186
rect 7658 8134 8832 8186
rect 1104 8112 8832 8134
rect 4816 8044 6684 8072
rect 4816 8016 4844 8044
rect 4798 7964 4804 8016
rect 4856 7964 4862 8016
rect 6546 7964 6552 8016
rect 6604 7964 6610 8016
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 4028 7908 5181 7936
rect 4028 7896 4034 7908
rect 5169 7905 5181 7908
rect 5215 7936 5227 7939
rect 6564 7936 6592 7964
rect 5215 7908 6592 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4663 7840 4844 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4154 7760 4160 7812
rect 4212 7800 4218 7812
rect 4709 7803 4767 7809
rect 4709 7800 4721 7803
rect 4212 7772 4721 7800
rect 4212 7760 4218 7772
rect 4709 7769 4721 7772
rect 4755 7769 4767 7803
rect 4709 7763 4767 7769
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 4816 7732 4844 7840
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 6656 7868 6684 8044
rect 7926 8032 7932 8084
rect 7984 8032 7990 8084
rect 7944 8004 7972 8032
rect 7944 7976 8340 8004
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 6963 7908 7573 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8312 7945 8340 7976
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 7892 7908 8217 7936
rect 7892 7896 7898 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 7190 7868 7196 7880
rect 6578 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7868 7254 7880
rect 7374 7868 7380 7880
rect 7248 7840 7380 7868
rect 7248 7828 7254 7840
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7800 7840 8125 7868
rect 7800 7828 7806 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 5350 7800 5356 7812
rect 4939 7772 5356 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 5718 7800 5724 7812
rect 5491 7772 5724 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 6972 7772 7972 7800
rect 6972 7760 6978 7772
rect 7944 7744 7972 7772
rect 5534 7732 5540 7744
rect 4816 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 7006 7692 7012 7744
rect 7064 7692 7070 7744
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 7926 7692 7932 7744
rect 7984 7692 7990 7744
rect 1104 7642 8832 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 8010 7642
rect 8062 7590 8074 7642
rect 8126 7590 8138 7642
rect 8190 7590 8202 7642
rect 8254 7590 8266 7642
rect 8318 7590 8832 7642
rect 1104 7568 8832 7590
rect 4154 7488 4160 7540
rect 4212 7488 4218 7540
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 5905 7531 5963 7537
rect 5905 7528 5917 7531
rect 5776 7500 5917 7528
rect 5776 7488 5782 7500
rect 5905 7497 5917 7500
rect 5951 7497 5963 7531
rect 7742 7528 7748 7540
rect 5905 7491 5963 7497
rect 6380 7500 7748 7528
rect 4172 7460 4200 7488
rect 3712 7432 4200 7460
rect 4249 7463 4307 7469
rect 3712 7401 3740 7432
rect 4249 7429 4261 7463
rect 4295 7460 4307 7463
rect 4448 7460 4476 7488
rect 4295 7432 4476 7460
rect 4295 7429 4307 7432
rect 4249 7423 4307 7429
rect 4798 7420 4804 7472
rect 4856 7420 4862 7472
rect 6380 7401 6408 7500
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 7374 7420 7380 7472
rect 7432 7420 7438 7472
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 5994 7324 6000 7336
rect 5767 7296 6000 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 3878 7148 3884 7200
rect 3936 7148 3942 7200
rect 6104 7188 6132 7355
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6604 7364 6653 7392
rect 6604 7352 6610 7364
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6564 7296 6929 7324
rect 6564 7265 6592 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 6549 7259 6607 7265
rect 6549 7225 6561 7259
rect 6595 7225 6607 7259
rect 6549 7219 6607 7225
rect 6914 7188 6920 7200
rect 6104 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 1104 7098 8832 7120
rect 1104 7046 2350 7098
rect 2402 7046 2414 7098
rect 2466 7046 2478 7098
rect 2530 7046 2542 7098
rect 2594 7046 2606 7098
rect 2658 7046 7350 7098
rect 7402 7046 7414 7098
rect 7466 7046 7478 7098
rect 7530 7046 7542 7098
rect 7594 7046 7606 7098
rect 7658 7046 8832 7098
rect 1104 7024 8832 7046
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 4046 6987 4104 6993
rect 4046 6984 4058 6987
rect 3936 6956 4058 6984
rect 3936 6944 3942 6956
rect 4046 6953 4058 6956
rect 4092 6953 4104 6987
rect 4046 6947 4104 6953
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5997 6987 6055 6993
rect 5997 6984 6009 6987
rect 5592 6956 6009 6984
rect 5592 6944 5598 6956
rect 5997 6953 6009 6956
rect 6043 6953 6055 6987
rect 5997 6947 6055 6953
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7745 6987 7803 6993
rect 7745 6984 7757 6987
rect 6972 6956 7757 6984
rect 6972 6944 6978 6956
rect 7745 6953 7757 6956
rect 7791 6953 7803 6987
rect 7745 6947 7803 6953
rect 6181 6919 6239 6925
rect 6181 6885 6193 6919
rect 6227 6885 6239 6919
rect 6181 6879 6239 6885
rect 6196 6848 6224 6879
rect 7006 6876 7012 6928
rect 7064 6876 7070 6928
rect 7024 6848 7052 6876
rect 6196 6820 7052 6848
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 7834 6848 7840 6860
rect 7607 6820 7840 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3804 6712 3832 6743
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 7285 6783 7343 6789
rect 7285 6780 7297 6783
rect 7156 6752 7297 6780
rect 7156 6740 7162 6752
rect 7285 6749 7297 6752
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 3970 6712 3976 6724
rect 3804 6684 3976 6712
rect 3970 6672 3976 6684
rect 4028 6672 4034 6724
rect 4798 6672 4804 6724
rect 4856 6672 4862 6724
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 6457 6715 6515 6721
rect 6457 6712 6469 6715
rect 5684 6684 6469 6712
rect 5684 6672 5690 6684
rect 6457 6681 6469 6684
rect 6503 6712 6515 6715
rect 7576 6712 7604 6811
rect 7834 6808 7840 6820
rect 7892 6848 7898 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 7892 6820 8309 6848
rect 7892 6808 7898 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 6503 6684 7604 6712
rect 6503 6681 6515 6684
rect 6457 6675 6515 6681
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 7834 6604 7840 6656
rect 7892 6644 7898 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 7892 6616 8125 6644
rect 7892 6604 7898 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 8205 6647 8263 6653
rect 8205 6613 8217 6647
rect 8251 6644 8263 6647
rect 8478 6644 8484 6656
rect 8251 6616 8484 6644
rect 8251 6613 8263 6616
rect 8205 6607 8263 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 1104 6554 8832 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 8010 6554
rect 8062 6502 8074 6554
rect 8126 6502 8138 6554
rect 8190 6502 8202 6554
rect 8254 6502 8266 6554
rect 8318 6502 8832 6554
rect 1104 6480 8832 6502
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7377 6443 7435 6449
rect 7377 6440 7389 6443
rect 7156 6412 7389 6440
rect 7156 6400 7162 6412
rect 7377 6409 7389 6412
rect 7423 6409 7435 6443
rect 7377 6403 7435 6409
rect 7834 6400 7840 6452
rect 7892 6400 7898 6452
rect 7650 6332 7656 6384
rect 7708 6332 7714 6384
rect 8386 6264 8392 6316
rect 8444 6264 8450 6316
rect 1104 6010 8832 6032
rect 1104 5958 2350 6010
rect 2402 5958 2414 6010
rect 2466 5958 2478 6010
rect 2530 5958 2542 6010
rect 2594 5958 2606 6010
rect 2658 5958 7350 6010
rect 7402 5958 7414 6010
rect 7466 5958 7478 6010
rect 7530 5958 7542 6010
rect 7594 5958 7606 6010
rect 7658 5958 8832 6010
rect 1104 5936 8832 5958
rect 8297 5899 8355 5905
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 8478 5896 8484 5908
rect 8343 5868 8484 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8846 5692 8852 5704
rect 8527 5664 8852 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 1104 5466 8832 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 8010 5466
rect 8062 5414 8074 5466
rect 8126 5414 8138 5466
rect 8190 5414 8202 5466
rect 8254 5414 8266 5466
rect 8318 5414 8832 5466
rect 1104 5392 8832 5414
rect 1104 4922 8832 4944
rect 1104 4870 2350 4922
rect 2402 4870 2414 4922
rect 2466 4870 2478 4922
rect 2530 4870 2542 4922
rect 2594 4870 2606 4922
rect 2658 4870 7350 4922
rect 7402 4870 7414 4922
rect 7466 4870 7478 4922
rect 7530 4870 7542 4922
rect 7594 4870 7606 4922
rect 7658 4870 8832 4922
rect 1104 4848 8832 4870
rect 1104 4378 8832 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 8010 4378
rect 8062 4326 8074 4378
rect 8126 4326 8138 4378
rect 8190 4326 8202 4378
rect 8254 4326 8266 4378
rect 8318 4326 8832 4378
rect 1104 4304 8832 4326
rect 1104 3834 8832 3856
rect 1104 3782 2350 3834
rect 2402 3782 2414 3834
rect 2466 3782 2478 3834
rect 2530 3782 2542 3834
rect 2594 3782 2606 3834
rect 2658 3782 7350 3834
rect 7402 3782 7414 3834
rect 7466 3782 7478 3834
rect 7530 3782 7542 3834
rect 7594 3782 7606 3834
rect 7658 3782 8832 3834
rect 1104 3760 8832 3782
rect 1104 3290 8832 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 8010 3290
rect 8062 3238 8074 3290
rect 8126 3238 8138 3290
rect 8190 3238 8202 3290
rect 8254 3238 8266 3290
rect 8318 3238 8832 3290
rect 1104 3216 8832 3238
rect 1854 3000 1860 3052
rect 1912 3000 1918 3052
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 2363 3012 2421 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 842 2796 848 2848
rect 900 2836 906 2848
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 900 2808 1685 2836
rect 900 2796 906 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 2130 2796 2136 2848
rect 2188 2796 2194 2848
rect 1104 2746 8832 2768
rect 1104 2694 2350 2746
rect 2402 2694 2414 2746
rect 2466 2694 2478 2746
rect 2530 2694 2542 2746
rect 2594 2694 2606 2746
rect 2658 2694 7350 2746
rect 7402 2694 7414 2746
rect 7466 2694 7478 2746
rect 7530 2694 7542 2746
rect 7594 2694 7606 2746
rect 7658 2694 8832 2746
rect 1104 2672 8832 2694
rect 7561 2635 7619 2641
rect 7561 2601 7573 2635
rect 7607 2632 7619 2635
rect 7742 2632 7748 2644
rect 7607 2604 7748 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 7926 2592 7932 2644
rect 7984 2592 7990 2644
rect 1854 2456 1860 2508
rect 1912 2456 1918 2508
rect 6638 2456 6644 2508
rect 6696 2456 6702 2508
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 5534 2428 5540 2440
rect 4479 2400 5540 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5868 2400 6377 2428
rect 5868 2388 5874 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 7944 2428 7972 2592
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7944 2400 8125 2428
rect 6365 2391 6423 2397
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 7650 2320 7656 2372
rect 7708 2320 7714 2372
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 9122 2360 9128 2372
rect 8527 2332 9128 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 4154 2252 4160 2304
rect 4212 2252 4218 2304
rect 1104 2202 8832 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 8010 2202
rect 8062 2150 8074 2202
rect 8126 2150 8138 2202
rect 8190 2150 8202 2202
rect 8254 2150 8266 2202
rect 8318 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 2350 77766 2402 77818
rect 2414 77766 2466 77818
rect 2478 77766 2530 77818
rect 2542 77766 2594 77818
rect 2606 77766 2658 77818
rect 7350 77766 7402 77818
rect 7414 77766 7466 77818
rect 7478 77766 7530 77818
rect 7542 77766 7594 77818
rect 7606 77766 7658 77818
rect 2688 77503 2740 77512
rect 2688 77469 2697 77503
rect 2697 77469 2731 77503
rect 2731 77469 2740 77503
rect 2688 77460 2740 77469
rect 5540 77392 5592 77444
rect 3010 77222 3062 77274
rect 3074 77222 3126 77274
rect 3138 77222 3190 77274
rect 3202 77222 3254 77274
rect 3266 77222 3318 77274
rect 8010 77222 8062 77274
rect 8074 77222 8126 77274
rect 8138 77222 8190 77274
rect 8202 77222 8254 77274
rect 8266 77222 8318 77274
rect 2350 76678 2402 76730
rect 2414 76678 2466 76730
rect 2478 76678 2530 76730
rect 2542 76678 2594 76730
rect 2606 76678 2658 76730
rect 7350 76678 7402 76730
rect 7414 76678 7466 76730
rect 7478 76678 7530 76730
rect 7542 76678 7594 76730
rect 7606 76678 7658 76730
rect 3010 76134 3062 76186
rect 3074 76134 3126 76186
rect 3138 76134 3190 76186
rect 3202 76134 3254 76186
rect 3266 76134 3318 76186
rect 8010 76134 8062 76186
rect 8074 76134 8126 76186
rect 8138 76134 8190 76186
rect 8202 76134 8254 76186
rect 8266 76134 8318 76186
rect 2350 75590 2402 75642
rect 2414 75590 2466 75642
rect 2478 75590 2530 75642
rect 2542 75590 2594 75642
rect 2606 75590 2658 75642
rect 7350 75590 7402 75642
rect 7414 75590 7466 75642
rect 7478 75590 7530 75642
rect 7542 75590 7594 75642
rect 7606 75590 7658 75642
rect 3010 75046 3062 75098
rect 3074 75046 3126 75098
rect 3138 75046 3190 75098
rect 3202 75046 3254 75098
rect 3266 75046 3318 75098
rect 8010 75046 8062 75098
rect 8074 75046 8126 75098
rect 8138 75046 8190 75098
rect 8202 75046 8254 75098
rect 8266 75046 8318 75098
rect 2350 74502 2402 74554
rect 2414 74502 2466 74554
rect 2478 74502 2530 74554
rect 2542 74502 2594 74554
rect 2606 74502 2658 74554
rect 7350 74502 7402 74554
rect 7414 74502 7466 74554
rect 7478 74502 7530 74554
rect 7542 74502 7594 74554
rect 7606 74502 7658 74554
rect 7932 74196 7984 74248
rect 8392 74103 8444 74112
rect 8392 74069 8401 74103
rect 8401 74069 8435 74103
rect 8435 74069 8444 74103
rect 8392 74060 8444 74069
rect 3010 73958 3062 74010
rect 3074 73958 3126 74010
rect 3138 73958 3190 74010
rect 3202 73958 3254 74010
rect 3266 73958 3318 74010
rect 8010 73958 8062 74010
rect 8074 73958 8126 74010
rect 8138 73958 8190 74010
rect 8202 73958 8254 74010
rect 8266 73958 8318 74010
rect 7748 73788 7800 73840
rect 5540 73720 5592 73772
rect 6368 73763 6420 73772
rect 6368 73729 6377 73763
rect 6377 73729 6411 73763
rect 6411 73729 6420 73763
rect 6368 73720 6420 73729
rect 6736 73695 6788 73704
rect 6736 73661 6745 73695
rect 6745 73661 6779 73695
rect 6779 73661 6788 73695
rect 6736 73652 6788 73661
rect 7012 73695 7064 73704
rect 7012 73661 7021 73695
rect 7021 73661 7055 73695
rect 7055 73661 7064 73695
rect 7012 73652 7064 73661
rect 6644 73516 6696 73568
rect 8024 73516 8076 73568
rect 2350 73414 2402 73466
rect 2414 73414 2466 73466
rect 2478 73414 2530 73466
rect 2542 73414 2594 73466
rect 2606 73414 2658 73466
rect 7350 73414 7402 73466
rect 7414 73414 7466 73466
rect 7478 73414 7530 73466
rect 7542 73414 7594 73466
rect 7606 73414 7658 73466
rect 7012 73312 7064 73364
rect 7840 73244 7892 73296
rect 5080 73151 5132 73160
rect 5080 73117 5089 73151
rect 5089 73117 5123 73151
rect 5123 73117 5132 73151
rect 5080 73108 5132 73117
rect 8024 73176 8076 73228
rect 5356 73083 5408 73092
rect 5356 73049 5365 73083
rect 5365 73049 5399 73083
rect 5399 73049 5408 73083
rect 5356 73040 5408 73049
rect 6644 73040 6696 73092
rect 6828 73015 6880 73024
rect 6828 72981 6837 73015
rect 6837 72981 6871 73015
rect 6871 72981 6880 73015
rect 6828 72972 6880 72981
rect 8024 73040 8076 73092
rect 7748 72972 7800 73024
rect 3010 72870 3062 72922
rect 3074 72870 3126 72922
rect 3138 72870 3190 72922
rect 3202 72870 3254 72922
rect 3266 72870 3318 72922
rect 8010 72870 8062 72922
rect 8074 72870 8126 72922
rect 8138 72870 8190 72922
rect 8202 72870 8254 72922
rect 8266 72870 8318 72922
rect 5356 72768 5408 72820
rect 6644 72768 6696 72820
rect 7932 72768 7984 72820
rect 6644 72632 6696 72684
rect 7012 72632 7064 72684
rect 6828 72607 6880 72616
rect 6828 72573 6837 72607
rect 6837 72573 6871 72607
rect 6871 72573 6880 72607
rect 6828 72564 6880 72573
rect 6460 72428 6512 72480
rect 7104 72428 7156 72480
rect 2350 72326 2402 72378
rect 2414 72326 2466 72378
rect 2478 72326 2530 72378
rect 2542 72326 2594 72378
rect 2606 72326 2658 72378
rect 7350 72326 7402 72378
rect 7414 72326 7466 72378
rect 7478 72326 7530 72378
rect 7542 72326 7594 72378
rect 7606 72326 7658 72378
rect 4436 72088 4488 72140
rect 5080 72088 5132 72140
rect 6736 72131 6788 72140
rect 6736 72097 6745 72131
rect 6745 72097 6779 72131
rect 6779 72097 6788 72131
rect 6736 72088 6788 72097
rect 7104 72088 7156 72140
rect 5080 71995 5132 72004
rect 5080 71961 5089 71995
rect 5089 71961 5123 71995
rect 5123 71961 5132 71995
rect 5080 71952 5132 71961
rect 5816 71884 5868 71936
rect 6552 72020 6604 72072
rect 7104 71952 7156 72004
rect 6552 71927 6604 71936
rect 6552 71893 6561 71927
rect 6561 71893 6595 71927
rect 6595 71893 6604 71927
rect 6552 71884 6604 71893
rect 7748 71884 7800 71936
rect 7932 71884 7984 71936
rect 3010 71782 3062 71834
rect 3074 71782 3126 71834
rect 3138 71782 3190 71834
rect 3202 71782 3254 71834
rect 3266 71782 3318 71834
rect 8010 71782 8062 71834
rect 8074 71782 8126 71834
rect 8138 71782 8190 71834
rect 8202 71782 8254 71834
rect 8266 71782 8318 71834
rect 5080 71680 5132 71732
rect 6828 71680 6880 71732
rect 7012 71680 7064 71732
rect 8484 71680 8536 71732
rect 7932 71612 7984 71664
rect 5908 71476 5960 71528
rect 6552 71476 6604 71528
rect 6460 71408 6512 71460
rect 7840 71519 7892 71528
rect 7840 71485 7849 71519
rect 7849 71485 7883 71519
rect 7883 71485 7892 71519
rect 7840 71476 7892 71485
rect 6092 71340 6144 71392
rect 2350 71238 2402 71290
rect 2414 71238 2466 71290
rect 2478 71238 2530 71290
rect 2542 71238 2594 71290
rect 2606 71238 2658 71290
rect 7350 71238 7402 71290
rect 7414 71238 7466 71290
rect 7478 71238 7530 71290
rect 7542 71238 7594 71290
rect 7606 71238 7658 71290
rect 6092 71043 6144 71052
rect 6092 71009 6101 71043
rect 6101 71009 6135 71043
rect 6135 71009 6144 71043
rect 6092 71000 6144 71009
rect 4988 70796 5040 70848
rect 5908 70975 5960 70984
rect 5908 70941 5917 70975
rect 5917 70941 5951 70975
rect 5951 70941 5960 70975
rect 5908 70932 5960 70941
rect 6920 70932 6972 70984
rect 7932 70932 7984 70984
rect 6184 70796 6236 70848
rect 7012 70839 7064 70848
rect 7012 70805 7021 70839
rect 7021 70805 7055 70839
rect 7055 70805 7064 70839
rect 7012 70796 7064 70805
rect 8392 70839 8444 70848
rect 8392 70805 8401 70839
rect 8401 70805 8435 70839
rect 8435 70805 8444 70839
rect 8392 70796 8444 70805
rect 3010 70694 3062 70746
rect 3074 70694 3126 70746
rect 3138 70694 3190 70746
rect 3202 70694 3254 70746
rect 3266 70694 3318 70746
rect 8010 70694 8062 70746
rect 8074 70694 8126 70746
rect 8138 70694 8190 70746
rect 8202 70694 8254 70746
rect 8266 70694 8318 70746
rect 4988 70524 5040 70576
rect 7012 70567 7064 70576
rect 7012 70533 7021 70567
rect 7021 70533 7055 70567
rect 7055 70533 7064 70567
rect 7012 70524 7064 70533
rect 7104 70524 7156 70576
rect 4436 70499 4488 70508
rect 4436 70465 4445 70499
rect 4445 70465 4479 70499
rect 4479 70465 4488 70499
rect 4436 70456 4488 70465
rect 5816 70456 5868 70508
rect 6184 70431 6236 70440
rect 6184 70397 6193 70431
rect 6193 70397 6227 70431
rect 6227 70397 6236 70431
rect 6184 70388 6236 70397
rect 6736 70499 6788 70508
rect 6736 70465 6745 70499
rect 6745 70465 6779 70499
rect 6779 70465 6788 70499
rect 6736 70456 6788 70465
rect 7012 70388 7064 70440
rect 8024 70320 8076 70372
rect 2350 70150 2402 70202
rect 2414 70150 2466 70202
rect 2478 70150 2530 70202
rect 2542 70150 2594 70202
rect 2606 70150 2658 70202
rect 7350 70150 7402 70202
rect 7414 70150 7466 70202
rect 7478 70150 7530 70202
rect 7542 70150 7594 70202
rect 7606 70150 7658 70202
rect 6920 70091 6972 70100
rect 6920 70057 6929 70091
rect 6929 70057 6963 70091
rect 6963 70057 6972 70091
rect 6920 70048 6972 70057
rect 7840 69912 7892 69964
rect 7932 69844 7984 69896
rect 5908 69708 5960 69760
rect 6184 69708 6236 69760
rect 3010 69606 3062 69658
rect 3074 69606 3126 69658
rect 3138 69606 3190 69658
rect 3202 69606 3254 69658
rect 3266 69606 3318 69658
rect 8010 69606 8062 69658
rect 8074 69606 8126 69658
rect 8138 69606 8190 69658
rect 8202 69606 8254 69658
rect 8266 69606 8318 69658
rect 4436 69411 4488 69420
rect 4436 69377 4445 69411
rect 4445 69377 4479 69411
rect 4479 69377 4488 69411
rect 4436 69368 4488 69377
rect 7104 69368 7156 69420
rect 8484 69368 8536 69420
rect 4712 69343 4764 69352
rect 4712 69309 4721 69343
rect 4721 69309 4755 69343
rect 4755 69309 4764 69343
rect 4712 69300 4764 69309
rect 6000 69300 6052 69352
rect 7840 69300 7892 69352
rect 6644 69164 6696 69216
rect 8392 69207 8444 69216
rect 8392 69173 8401 69207
rect 8401 69173 8435 69207
rect 8435 69173 8444 69207
rect 8392 69164 8444 69173
rect 2350 69062 2402 69114
rect 2414 69062 2466 69114
rect 2478 69062 2530 69114
rect 2542 69062 2594 69114
rect 2606 69062 2658 69114
rect 7350 69062 7402 69114
rect 7414 69062 7466 69114
rect 7478 69062 7530 69114
rect 7542 69062 7594 69114
rect 7606 69062 7658 69114
rect 4712 68960 4764 69012
rect 8484 69003 8536 69012
rect 8484 68969 8493 69003
rect 8493 68969 8527 69003
rect 8527 68969 8536 69003
rect 8484 68960 8536 68969
rect 6000 68867 6052 68876
rect 6000 68833 6009 68867
rect 6009 68833 6043 68867
rect 6043 68833 6052 68867
rect 6000 68824 6052 68833
rect 6276 68824 6328 68876
rect 5908 68799 5960 68808
rect 5908 68765 5917 68799
rect 5917 68765 5951 68799
rect 5951 68765 5960 68799
rect 5908 68756 5960 68765
rect 6644 68756 6696 68808
rect 6736 68799 6788 68808
rect 6736 68765 6745 68799
rect 6745 68765 6779 68799
rect 6779 68765 6788 68799
rect 6736 68756 6788 68765
rect 7104 68688 7156 68740
rect 3010 68518 3062 68570
rect 3074 68518 3126 68570
rect 3138 68518 3190 68570
rect 3202 68518 3254 68570
rect 3266 68518 3318 68570
rect 8010 68518 8062 68570
rect 8074 68518 8126 68570
rect 8138 68518 8190 68570
rect 8202 68518 8254 68570
rect 8266 68518 8318 68570
rect 6000 68416 6052 68468
rect 6552 68280 6604 68332
rect 6828 68212 6880 68264
rect 7840 68212 7892 68264
rect 5172 68119 5224 68128
rect 5172 68085 5181 68119
rect 5181 68085 5215 68119
rect 5215 68085 5224 68119
rect 5172 68076 5224 68085
rect 7748 68076 7800 68128
rect 8392 68119 8444 68128
rect 8392 68085 8401 68119
rect 8401 68085 8435 68119
rect 8435 68085 8444 68119
rect 8392 68076 8444 68085
rect 2350 67974 2402 68026
rect 2414 67974 2466 68026
rect 2478 67974 2530 68026
rect 2542 67974 2594 68026
rect 2606 67974 2658 68026
rect 7350 67974 7402 68026
rect 7414 67974 7466 68026
rect 7478 67974 7530 68026
rect 7542 67974 7594 68026
rect 7606 67974 7658 68026
rect 6552 67915 6604 67924
rect 6552 67881 6561 67915
rect 6561 67881 6595 67915
rect 6595 67881 6604 67915
rect 6552 67872 6604 67881
rect 4436 67736 4488 67788
rect 5172 67736 5224 67788
rect 7012 67736 7064 67788
rect 7656 67736 7708 67788
rect 6736 67711 6788 67720
rect 6736 67677 6745 67711
rect 6745 67677 6779 67711
rect 6779 67677 6788 67711
rect 6736 67668 6788 67677
rect 6092 67532 6144 67584
rect 7012 67643 7064 67652
rect 7012 67609 7021 67643
rect 7021 67609 7055 67643
rect 7055 67609 7064 67643
rect 7012 67600 7064 67609
rect 7104 67600 7156 67652
rect 3010 67430 3062 67482
rect 3074 67430 3126 67482
rect 3138 67430 3190 67482
rect 3202 67430 3254 67482
rect 3266 67430 3318 67482
rect 8010 67430 8062 67482
rect 8074 67430 8126 67482
rect 8138 67430 8190 67482
rect 8202 67430 8254 67482
rect 8266 67430 8318 67482
rect 6552 67328 6604 67380
rect 7012 67328 7064 67380
rect 7748 67328 7800 67380
rect 6920 67260 6972 67312
rect 8484 67192 8536 67244
rect 6828 67124 6880 67176
rect 6368 67031 6420 67040
rect 6368 66997 6377 67031
rect 6377 66997 6411 67031
rect 6411 66997 6420 67031
rect 6368 66988 6420 66997
rect 8392 67031 8444 67040
rect 8392 66997 8401 67031
rect 8401 66997 8435 67031
rect 8435 66997 8444 67031
rect 8392 66988 8444 66997
rect 2350 66886 2402 66938
rect 2414 66886 2466 66938
rect 2478 66886 2530 66938
rect 2542 66886 2594 66938
rect 2606 66886 2658 66938
rect 7350 66886 7402 66938
rect 7414 66886 7466 66938
rect 7478 66886 7530 66938
rect 7542 66886 7594 66938
rect 7606 66886 7658 66938
rect 6920 66784 6972 66836
rect 4436 66648 4488 66700
rect 6092 66580 6144 66632
rect 7012 66580 7064 66632
rect 7104 66580 7156 66632
rect 7840 66580 7892 66632
rect 5080 66555 5132 66564
rect 5080 66521 5089 66555
rect 5089 66521 5123 66555
rect 5123 66521 5132 66555
rect 5080 66512 5132 66521
rect 5724 66444 5776 66496
rect 6736 66512 6788 66564
rect 7656 66487 7708 66496
rect 7656 66453 7665 66487
rect 7665 66453 7699 66487
rect 7699 66453 7708 66487
rect 7656 66444 7708 66453
rect 8484 66444 8536 66496
rect 3010 66342 3062 66394
rect 3074 66342 3126 66394
rect 3138 66342 3190 66394
rect 3202 66342 3254 66394
rect 3266 66342 3318 66394
rect 8010 66342 8062 66394
rect 8074 66342 8126 66394
rect 8138 66342 8190 66394
rect 8202 66342 8254 66394
rect 8266 66342 8318 66394
rect 5080 66240 5132 66292
rect 6368 66240 6420 66292
rect 7656 66240 7708 66292
rect 8484 66283 8536 66292
rect 8484 66249 8493 66283
rect 8493 66249 8527 66283
rect 8527 66249 8536 66283
rect 8484 66240 8536 66249
rect 7012 66172 7064 66224
rect 6736 66079 6788 66088
rect 6736 66045 6745 66079
rect 6745 66045 6779 66079
rect 6779 66045 6788 66079
rect 6736 66036 6788 66045
rect 2350 65798 2402 65850
rect 2414 65798 2466 65850
rect 2478 65798 2530 65850
rect 2542 65798 2594 65850
rect 2606 65798 2658 65850
rect 7350 65798 7402 65850
rect 7414 65798 7466 65850
rect 7478 65798 7530 65850
rect 7542 65798 7594 65850
rect 7606 65798 7658 65850
rect 4436 65560 4488 65612
rect 5816 65560 5868 65612
rect 6828 65560 6880 65612
rect 6092 65492 6144 65544
rect 6920 65492 6972 65544
rect 7932 65492 7984 65544
rect 5080 65467 5132 65476
rect 5080 65433 5089 65467
rect 5089 65433 5123 65467
rect 5123 65433 5132 65467
rect 5080 65424 5132 65433
rect 6920 65399 6972 65408
rect 6920 65365 6929 65399
rect 6929 65365 6963 65399
rect 6963 65365 6972 65399
rect 6920 65356 6972 65365
rect 7748 65356 7800 65408
rect 8392 65399 8444 65408
rect 8392 65365 8401 65399
rect 8401 65365 8435 65399
rect 8435 65365 8444 65399
rect 8392 65356 8444 65365
rect 3010 65254 3062 65306
rect 3074 65254 3126 65306
rect 3138 65254 3190 65306
rect 3202 65254 3254 65306
rect 3266 65254 3318 65306
rect 8010 65254 8062 65306
rect 8074 65254 8126 65306
rect 8138 65254 8190 65306
rect 8202 65254 8254 65306
rect 8266 65254 8318 65306
rect 5080 65152 5132 65204
rect 6920 65152 6972 65204
rect 4436 65084 4488 65136
rect 5540 65059 5592 65068
rect 5540 65025 5549 65059
rect 5549 65025 5583 65059
rect 5583 65025 5592 65059
rect 5540 65016 5592 65025
rect 7840 65084 7892 65136
rect 7104 65016 7156 65068
rect 7012 64855 7064 64864
rect 7012 64821 7021 64855
rect 7021 64821 7055 64855
rect 7055 64821 7064 64855
rect 7012 64812 7064 64821
rect 8208 64855 8260 64864
rect 8208 64821 8217 64855
rect 8217 64821 8251 64855
rect 8251 64821 8260 64855
rect 8208 64812 8260 64821
rect 2350 64710 2402 64762
rect 2414 64710 2466 64762
rect 2478 64710 2530 64762
rect 2542 64710 2594 64762
rect 2606 64710 2658 64762
rect 7350 64710 7402 64762
rect 7414 64710 7466 64762
rect 7478 64710 7530 64762
rect 7542 64710 7594 64762
rect 7606 64710 7658 64762
rect 7012 64515 7064 64524
rect 7012 64481 7021 64515
rect 7021 64481 7055 64515
rect 7055 64481 7064 64515
rect 7012 64472 7064 64481
rect 7656 64472 7708 64524
rect 8208 64472 8260 64524
rect 6460 64447 6512 64456
rect 6460 64413 6469 64447
rect 6469 64413 6503 64447
rect 6503 64413 6512 64447
rect 6460 64404 6512 64413
rect 6736 64447 6788 64456
rect 6736 64413 6745 64447
rect 6745 64413 6779 64447
rect 6779 64413 6788 64447
rect 6736 64404 6788 64413
rect 6644 64311 6696 64320
rect 6644 64277 6653 64311
rect 6653 64277 6687 64311
rect 6687 64277 6696 64311
rect 6644 64268 6696 64277
rect 7932 64268 7984 64320
rect 3010 64166 3062 64218
rect 3074 64166 3126 64218
rect 3138 64166 3190 64218
rect 3202 64166 3254 64218
rect 3266 64166 3318 64218
rect 8010 64166 8062 64218
rect 8074 64166 8126 64218
rect 8138 64166 8190 64218
rect 8202 64166 8254 64218
rect 8266 64166 8318 64218
rect 6644 64064 6696 64116
rect 7012 64064 7064 64116
rect 7656 64064 7708 64116
rect 5908 63928 5960 63980
rect 5724 63903 5776 63912
rect 5724 63869 5733 63903
rect 5733 63869 5767 63903
rect 5767 63869 5776 63903
rect 5724 63860 5776 63869
rect 5816 63903 5868 63912
rect 5816 63869 5825 63903
rect 5825 63869 5859 63903
rect 5859 63869 5868 63903
rect 5816 63860 5868 63869
rect 4804 63767 4856 63776
rect 4804 63733 4813 63767
rect 4813 63733 4847 63767
rect 4847 63733 4856 63767
rect 4804 63724 4856 63733
rect 6736 63724 6788 63776
rect 8208 63767 8260 63776
rect 8208 63733 8217 63767
rect 8217 63733 8251 63767
rect 8251 63733 8260 63767
rect 8208 63724 8260 63733
rect 2350 63622 2402 63674
rect 2414 63622 2466 63674
rect 2478 63622 2530 63674
rect 2542 63622 2594 63674
rect 2606 63622 2658 63674
rect 7350 63622 7402 63674
rect 7414 63622 7466 63674
rect 7478 63622 7530 63674
rect 7542 63622 7594 63674
rect 7606 63622 7658 63674
rect 4804 63520 4856 63572
rect 5724 63520 5776 63572
rect 4344 63427 4396 63436
rect 4344 63393 4353 63427
rect 4353 63393 4387 63427
rect 4387 63393 4396 63427
rect 4344 63384 4396 63393
rect 6460 63520 6512 63572
rect 7840 63520 7892 63572
rect 7104 63452 7156 63504
rect 7288 63452 7340 63504
rect 8484 63520 8536 63572
rect 7840 63427 7892 63436
rect 7840 63393 7849 63427
rect 7849 63393 7883 63427
rect 7883 63393 7892 63427
rect 7840 63384 7892 63393
rect 5908 63248 5960 63300
rect 8208 63316 8260 63368
rect 7104 63248 7156 63300
rect 7288 63248 7340 63300
rect 7932 63248 7984 63300
rect 6644 63180 6696 63232
rect 3010 63078 3062 63130
rect 3074 63078 3126 63130
rect 3138 63078 3190 63130
rect 3202 63078 3254 63130
rect 3266 63078 3318 63130
rect 8010 63078 8062 63130
rect 8074 63078 8126 63130
rect 8138 63078 8190 63130
rect 8202 63078 8254 63130
rect 8266 63078 8318 63130
rect 5724 62976 5776 63028
rect 8024 62840 8076 62892
rect 5908 62772 5960 62824
rect 6092 62772 6144 62824
rect 4712 62636 4764 62688
rect 8392 62679 8444 62688
rect 8392 62645 8401 62679
rect 8401 62645 8435 62679
rect 8435 62645 8444 62679
rect 8392 62636 8444 62645
rect 2350 62534 2402 62586
rect 2414 62534 2466 62586
rect 2478 62534 2530 62586
rect 2542 62534 2594 62586
rect 2606 62534 2658 62586
rect 7350 62534 7402 62586
rect 7414 62534 7466 62586
rect 7478 62534 7530 62586
rect 7542 62534 7594 62586
rect 7606 62534 7658 62586
rect 4344 62339 4396 62348
rect 4344 62305 4353 62339
rect 4353 62305 4387 62339
rect 4387 62305 4396 62339
rect 4344 62296 4396 62305
rect 4712 62296 4764 62348
rect 7104 62432 7156 62484
rect 7012 62296 7064 62348
rect 6460 62271 6512 62280
rect 6460 62237 6469 62271
rect 6469 62237 6503 62271
rect 6503 62237 6512 62271
rect 6460 62228 6512 62237
rect 6736 62271 6788 62280
rect 6736 62237 6745 62271
rect 6745 62237 6779 62271
rect 6779 62237 6788 62271
rect 6736 62228 6788 62237
rect 6092 62135 6144 62144
rect 6092 62101 6101 62135
rect 6101 62101 6135 62135
rect 6135 62101 6144 62135
rect 6092 62092 6144 62101
rect 7104 62092 7156 62144
rect 8024 62092 8076 62144
rect 3010 61990 3062 62042
rect 3074 61990 3126 62042
rect 3138 61990 3190 62042
rect 3202 61990 3254 62042
rect 3266 61990 3318 62042
rect 8010 61990 8062 62042
rect 8074 61990 8126 62042
rect 8138 61990 8190 62042
rect 8202 61990 8254 62042
rect 8266 61990 8318 62042
rect 6460 61888 6512 61940
rect 7104 61931 7156 61940
rect 7104 61897 7113 61931
rect 7113 61897 7147 61931
rect 7147 61897 7156 61931
rect 7104 61888 7156 61897
rect 6092 61820 6144 61872
rect 7104 61548 7156 61600
rect 2350 61446 2402 61498
rect 2414 61446 2466 61498
rect 2478 61446 2530 61498
rect 2542 61446 2594 61498
rect 2606 61446 2658 61498
rect 7350 61446 7402 61498
rect 7414 61446 7466 61498
rect 7478 61446 7530 61498
rect 7542 61446 7594 61498
rect 7606 61446 7658 61498
rect 4344 61208 4396 61260
rect 6828 61183 6880 61192
rect 6828 61149 6837 61183
rect 6837 61149 6871 61183
rect 6871 61149 6880 61183
rect 6828 61140 6880 61149
rect 7748 61140 7800 61192
rect 4712 61115 4764 61124
rect 4712 61081 4721 61115
rect 4721 61081 4755 61115
rect 4755 61081 4764 61115
rect 4712 61072 4764 61081
rect 6920 61072 6972 61124
rect 7932 61072 7984 61124
rect 5724 61004 5776 61056
rect 7012 61047 7064 61056
rect 7012 61013 7021 61047
rect 7021 61013 7055 61047
rect 7055 61013 7064 61047
rect 7012 61004 7064 61013
rect 7104 61004 7156 61056
rect 7380 61047 7432 61056
rect 7380 61013 7389 61047
rect 7389 61013 7423 61047
rect 7423 61013 7432 61047
rect 7380 61004 7432 61013
rect 8392 61047 8444 61056
rect 8392 61013 8401 61047
rect 8401 61013 8435 61047
rect 8435 61013 8444 61047
rect 8392 61004 8444 61013
rect 3010 60902 3062 60954
rect 3074 60902 3126 60954
rect 3138 60902 3190 60954
rect 3202 60902 3254 60954
rect 3266 60902 3318 60954
rect 8010 60902 8062 60954
rect 8074 60902 8126 60954
rect 8138 60902 8190 60954
rect 8202 60902 8254 60954
rect 8266 60902 8318 60954
rect 4712 60800 4764 60852
rect 6092 60800 6144 60852
rect 7104 60800 7156 60852
rect 6920 60732 6972 60784
rect 7012 60775 7064 60784
rect 7012 60741 7021 60775
rect 7021 60741 7055 60775
rect 7055 60741 7064 60775
rect 7012 60732 7064 60741
rect 7380 60800 7432 60852
rect 8024 60800 8076 60852
rect 5632 60707 5684 60716
rect 5632 60673 5641 60707
rect 5641 60673 5675 60707
rect 5675 60673 5684 60707
rect 5632 60664 5684 60673
rect 5908 60596 5960 60648
rect 6736 60639 6788 60648
rect 6736 60605 6745 60639
rect 6745 60605 6779 60639
rect 6779 60605 6788 60639
rect 6736 60596 6788 60605
rect 7012 60596 7064 60648
rect 7380 60596 7432 60648
rect 7012 60460 7064 60512
rect 7748 60460 7800 60512
rect 2350 60358 2402 60410
rect 2414 60358 2466 60410
rect 2478 60358 2530 60410
rect 2542 60358 2594 60410
rect 2606 60358 2658 60410
rect 7350 60358 7402 60410
rect 7414 60358 7466 60410
rect 7478 60358 7530 60410
rect 7542 60358 7594 60410
rect 7606 60358 7658 60410
rect 6828 60256 6880 60308
rect 5908 60120 5960 60172
rect 7012 60095 7064 60104
rect 7012 60061 7021 60095
rect 7021 60061 7055 60095
rect 7055 60061 7064 60095
rect 7012 60052 7064 60061
rect 5724 59984 5776 60036
rect 4896 59959 4948 59968
rect 4896 59925 4905 59959
rect 4905 59925 4939 59959
rect 4939 59925 4948 59959
rect 4896 59916 4948 59925
rect 6184 59916 6236 59968
rect 7012 59916 7064 59968
rect 8024 60120 8076 60172
rect 7748 60052 7800 60104
rect 8392 59959 8444 59968
rect 8392 59925 8401 59959
rect 8401 59925 8435 59959
rect 8435 59925 8444 59959
rect 8392 59916 8444 59925
rect 3010 59814 3062 59866
rect 3074 59814 3126 59866
rect 3138 59814 3190 59866
rect 3202 59814 3254 59866
rect 3266 59814 3318 59866
rect 8010 59814 8062 59866
rect 8074 59814 8126 59866
rect 8138 59814 8190 59866
rect 8202 59814 8254 59866
rect 8266 59814 8318 59866
rect 4896 59712 4948 59764
rect 4436 59619 4488 59628
rect 4436 59585 4445 59619
rect 4445 59585 4479 59619
rect 4479 59585 4488 59619
rect 4436 59576 4488 59585
rect 6460 59619 6512 59628
rect 6460 59585 6469 59619
rect 6469 59585 6503 59619
rect 6503 59585 6512 59619
rect 6460 59576 6512 59585
rect 6736 59551 6788 59560
rect 6736 59517 6745 59551
rect 6745 59517 6779 59551
rect 6779 59517 6788 59551
rect 6736 59508 6788 59517
rect 7104 59508 7156 59560
rect 5724 59372 5776 59424
rect 6184 59415 6236 59424
rect 6184 59381 6193 59415
rect 6193 59381 6227 59415
rect 6227 59381 6236 59415
rect 6184 59372 6236 59381
rect 7104 59372 7156 59424
rect 7748 59372 7800 59424
rect 2350 59270 2402 59322
rect 2414 59270 2466 59322
rect 2478 59270 2530 59322
rect 2542 59270 2594 59322
rect 2606 59270 2658 59322
rect 7350 59270 7402 59322
rect 7414 59270 7466 59322
rect 7478 59270 7530 59322
rect 7542 59270 7594 59322
rect 7606 59270 7658 59322
rect 6460 59168 6512 59220
rect 7012 59100 7064 59152
rect 5908 59075 5960 59084
rect 5908 59041 5917 59075
rect 5917 59041 5951 59075
rect 5951 59041 5960 59075
rect 5908 59032 5960 59041
rect 6184 59032 6236 59084
rect 7104 59007 7156 59016
rect 7104 58973 7113 59007
rect 7113 58973 7147 59007
rect 7147 58973 7156 59007
rect 7104 58964 7156 58973
rect 7748 58896 7800 58948
rect 5264 58871 5316 58880
rect 5264 58837 5273 58871
rect 5273 58837 5307 58871
rect 5307 58837 5316 58871
rect 5264 58828 5316 58837
rect 6000 58828 6052 58880
rect 8484 58828 8536 58880
rect 3010 58726 3062 58778
rect 3074 58726 3126 58778
rect 3138 58726 3190 58778
rect 3202 58726 3254 58778
rect 3266 58726 3318 58778
rect 8010 58726 8062 58778
rect 8074 58726 8126 58778
rect 8138 58726 8190 58778
rect 8202 58726 8254 58778
rect 8266 58726 8318 58778
rect 4712 58599 4764 58608
rect 4712 58565 4721 58599
rect 4721 58565 4755 58599
rect 4755 58565 4764 58599
rect 4712 58556 4764 58565
rect 5724 58488 5776 58540
rect 6460 58531 6512 58540
rect 6460 58497 6469 58531
rect 6469 58497 6503 58531
rect 6503 58497 6512 58531
rect 6460 58488 6512 58497
rect 6736 58463 6788 58472
rect 6736 58429 6745 58463
rect 6745 58429 6779 58463
rect 6779 58429 6788 58463
rect 6736 58420 6788 58429
rect 6000 58284 6052 58336
rect 7104 58284 7156 58336
rect 7748 58284 7800 58336
rect 2350 58182 2402 58234
rect 2414 58182 2466 58234
rect 2478 58182 2530 58234
rect 2542 58182 2594 58234
rect 2606 58182 2658 58234
rect 7350 58182 7402 58234
rect 7414 58182 7466 58234
rect 7478 58182 7530 58234
rect 7542 58182 7594 58234
rect 7606 58182 7658 58234
rect 4712 58080 4764 58132
rect 6460 58080 6512 58132
rect 7012 57944 7064 57996
rect 7748 57944 7800 57996
rect 5264 57876 5316 57928
rect 7104 57919 7156 57928
rect 7104 57885 7113 57919
rect 7113 57885 7147 57919
rect 7147 57885 7156 57919
rect 7104 57876 7156 57885
rect 6460 57808 6512 57860
rect 6000 57740 6052 57792
rect 7656 57740 7708 57792
rect 3010 57638 3062 57690
rect 3074 57638 3126 57690
rect 3138 57638 3190 57690
rect 3202 57638 3254 57690
rect 3266 57638 3318 57690
rect 8010 57638 8062 57690
rect 8074 57638 8126 57690
rect 8138 57638 8190 57690
rect 8202 57638 8254 57690
rect 8266 57638 8318 57690
rect 5724 57468 5776 57520
rect 6828 57443 6880 57452
rect 6828 57409 6837 57443
rect 6837 57409 6871 57443
rect 6871 57409 6880 57443
rect 6828 57400 6880 57409
rect 7104 57400 7156 57452
rect 4712 57375 4764 57384
rect 4712 57341 4721 57375
rect 4721 57341 4755 57375
rect 4755 57341 4764 57375
rect 4712 57332 4764 57341
rect 7656 57332 7708 57384
rect 8024 57332 8076 57384
rect 6092 57196 6144 57248
rect 6184 57239 6236 57248
rect 6184 57205 6193 57239
rect 6193 57205 6227 57239
rect 6227 57205 6236 57239
rect 6184 57196 6236 57205
rect 7012 57239 7064 57248
rect 7012 57205 7021 57239
rect 7021 57205 7055 57239
rect 7055 57205 7064 57239
rect 7012 57196 7064 57205
rect 8576 57196 8628 57248
rect 2350 57094 2402 57146
rect 2414 57094 2466 57146
rect 2478 57094 2530 57146
rect 2542 57094 2594 57146
rect 2606 57094 2658 57146
rect 7350 57094 7402 57146
rect 7414 57094 7466 57146
rect 7478 57094 7530 57146
rect 7542 57094 7594 57146
rect 7606 57094 7658 57146
rect 4712 56992 4764 57044
rect 6276 56992 6328 57044
rect 5908 56856 5960 56908
rect 6092 56856 6144 56908
rect 6736 56899 6788 56908
rect 6736 56865 6745 56899
rect 6745 56865 6779 56899
rect 6779 56865 6788 56899
rect 6736 56856 6788 56865
rect 7012 56899 7064 56908
rect 7012 56865 7021 56899
rect 7021 56865 7055 56899
rect 7055 56865 7064 56899
rect 7012 56856 7064 56865
rect 7104 56856 7156 56908
rect 6000 56788 6052 56840
rect 6276 56788 6328 56840
rect 8024 56788 8076 56840
rect 5632 56652 5684 56704
rect 7656 56652 7708 56704
rect 3010 56550 3062 56602
rect 3074 56550 3126 56602
rect 3138 56550 3190 56602
rect 3202 56550 3254 56602
rect 3266 56550 3318 56602
rect 8010 56550 8062 56602
rect 8074 56550 8126 56602
rect 8138 56550 8190 56602
rect 8202 56550 8254 56602
rect 8266 56550 8318 56602
rect 6460 56448 6512 56500
rect 6828 56448 6880 56500
rect 7104 56491 7156 56500
rect 7104 56457 7113 56491
rect 7113 56457 7147 56491
rect 7147 56457 7156 56491
rect 7104 56448 7156 56457
rect 5632 56423 5684 56432
rect 5632 56389 5641 56423
rect 5641 56389 5675 56423
rect 5675 56389 5684 56423
rect 5632 56380 5684 56389
rect 6184 56380 6236 56432
rect 6368 56312 6420 56364
rect 5632 56244 5684 56296
rect 5908 56287 5960 56296
rect 5908 56253 5917 56287
rect 5917 56253 5951 56287
rect 5951 56253 5960 56287
rect 5908 56244 5960 56253
rect 6920 56244 6972 56296
rect 7748 56244 7800 56296
rect 6828 56176 6880 56228
rect 7932 56176 7984 56228
rect 4896 56108 4948 56160
rect 7656 56108 7708 56160
rect 8024 56108 8076 56160
rect 2350 56006 2402 56058
rect 2414 56006 2466 56058
rect 2478 56006 2530 56058
rect 2542 56006 2594 56058
rect 2606 56006 2658 56058
rect 7350 56006 7402 56058
rect 7414 56006 7466 56058
rect 7478 56006 7530 56058
rect 7542 56006 7594 56058
rect 7606 56006 7658 56058
rect 6460 55836 6512 55888
rect 4896 55768 4948 55820
rect 6736 55811 6788 55820
rect 6736 55777 6745 55811
rect 6745 55777 6779 55811
rect 6779 55777 6788 55811
rect 6736 55768 6788 55777
rect 4436 55700 4488 55752
rect 5908 55700 5960 55752
rect 6460 55743 6512 55752
rect 6460 55709 6469 55743
rect 6469 55709 6503 55743
rect 6503 55709 6512 55743
rect 6460 55700 6512 55709
rect 8024 55700 8076 55752
rect 5632 55564 5684 55616
rect 6276 55607 6328 55616
rect 6276 55573 6285 55607
rect 6285 55573 6319 55607
rect 6319 55573 6328 55607
rect 6276 55564 6328 55573
rect 8484 55607 8536 55616
rect 8484 55573 8493 55607
rect 8493 55573 8527 55607
rect 8527 55573 8536 55607
rect 8484 55564 8536 55573
rect 3010 55462 3062 55514
rect 3074 55462 3126 55514
rect 3138 55462 3190 55514
rect 3202 55462 3254 55514
rect 3266 55462 3318 55514
rect 8010 55462 8062 55514
rect 8074 55462 8126 55514
rect 8138 55462 8190 55514
rect 8202 55462 8254 55514
rect 8266 55462 8318 55514
rect 6276 55360 6328 55412
rect 6460 55360 6512 55412
rect 6276 55224 6328 55276
rect 6644 55224 6696 55276
rect 8484 55267 8536 55276
rect 8484 55233 8493 55267
rect 8493 55233 8527 55267
rect 8527 55233 8536 55267
rect 8484 55224 8536 55233
rect 6920 55156 6972 55208
rect 2350 54918 2402 54970
rect 2414 54918 2466 54970
rect 2478 54918 2530 54970
rect 2542 54918 2594 54970
rect 2606 54918 2658 54970
rect 7350 54918 7402 54970
rect 7414 54918 7466 54970
rect 7478 54918 7530 54970
rect 7542 54918 7594 54970
rect 7606 54918 7658 54970
rect 8208 54816 8260 54868
rect 7656 54748 7708 54800
rect 7932 54748 7984 54800
rect 4436 54612 4488 54664
rect 5908 54612 5960 54664
rect 7932 54612 7984 54664
rect 8484 54612 8536 54664
rect 4804 54587 4856 54596
rect 4804 54553 4813 54587
rect 4813 54553 4847 54587
rect 4847 54553 4856 54587
rect 4804 54544 4856 54553
rect 5816 54476 5868 54528
rect 8392 54519 8444 54528
rect 8392 54485 8401 54519
rect 8401 54485 8435 54519
rect 8435 54485 8444 54519
rect 8392 54476 8444 54485
rect 3010 54374 3062 54426
rect 3074 54374 3126 54426
rect 3138 54374 3190 54426
rect 3202 54374 3254 54426
rect 3266 54374 3318 54426
rect 8010 54374 8062 54426
rect 8074 54374 8126 54426
rect 8138 54374 8190 54426
rect 8202 54374 8254 54426
rect 8266 54374 8318 54426
rect 4804 54272 4856 54324
rect 5632 54315 5684 54324
rect 5632 54281 5641 54315
rect 5641 54281 5675 54315
rect 5675 54281 5684 54315
rect 5632 54272 5684 54281
rect 7656 54204 7708 54256
rect 6460 54179 6512 54188
rect 6460 54145 6469 54179
rect 6469 54145 6503 54179
rect 6503 54145 6512 54179
rect 6460 54136 6512 54145
rect 6736 54179 6788 54188
rect 6736 54145 6745 54179
rect 6745 54145 6779 54179
rect 6779 54145 6788 54179
rect 6736 54136 6788 54145
rect 6184 54068 6236 54120
rect 7656 54068 7708 54120
rect 8116 54000 8168 54052
rect 5816 53932 5868 53984
rect 7012 53932 7064 53984
rect 8024 53932 8076 53984
rect 2350 53830 2402 53882
rect 2414 53830 2466 53882
rect 2478 53830 2530 53882
rect 2542 53830 2594 53882
rect 2606 53830 2658 53882
rect 7350 53830 7402 53882
rect 7414 53830 7466 53882
rect 7478 53830 7530 53882
rect 7542 53830 7594 53882
rect 7606 53830 7658 53882
rect 6460 53728 6512 53780
rect 6184 53592 6236 53644
rect 6644 53592 6696 53644
rect 6920 53592 6972 53644
rect 4988 53431 5040 53440
rect 4988 53397 4997 53431
rect 4997 53397 5031 53431
rect 5031 53397 5040 53431
rect 4988 53388 5040 53397
rect 7012 53567 7064 53576
rect 7012 53533 7021 53567
rect 7021 53533 7055 53567
rect 7055 53533 7064 53567
rect 7012 53524 7064 53533
rect 5816 53456 5868 53508
rect 6184 53388 6236 53440
rect 3010 53286 3062 53338
rect 3074 53286 3126 53338
rect 3138 53286 3190 53338
rect 3202 53286 3254 53338
rect 3266 53286 3318 53338
rect 8010 53286 8062 53338
rect 8074 53286 8126 53338
rect 8138 53286 8190 53338
rect 8202 53286 8254 53338
rect 8266 53286 8318 53338
rect 4988 53184 5040 53236
rect 7932 53184 7984 53236
rect 6460 53091 6512 53100
rect 6460 53057 6469 53091
rect 6469 53057 6503 53091
rect 6503 53057 6512 53091
rect 6460 53048 6512 53057
rect 6736 53091 6788 53100
rect 6736 53057 6745 53091
rect 6745 53057 6779 53091
rect 6779 53057 6788 53091
rect 6736 53048 6788 53057
rect 4436 53023 4488 53032
rect 4436 52989 4445 53023
rect 4445 52989 4479 53023
rect 4479 52989 4488 53023
rect 4436 52980 4488 52989
rect 5908 52980 5960 53032
rect 6184 52887 6236 52896
rect 6184 52853 6193 52887
rect 6193 52853 6227 52887
rect 6227 52853 6236 52887
rect 6184 52844 6236 52853
rect 8208 52844 8260 52896
rect 2350 52742 2402 52794
rect 2414 52742 2466 52794
rect 2478 52742 2530 52794
rect 2542 52742 2594 52794
rect 2606 52742 2658 52794
rect 7350 52742 7402 52794
rect 7414 52742 7466 52794
rect 7478 52742 7530 52794
rect 7542 52742 7594 52794
rect 7606 52742 7658 52794
rect 6460 52640 6512 52692
rect 8392 52683 8444 52692
rect 8392 52649 8401 52683
rect 8401 52649 8435 52683
rect 8435 52649 8444 52683
rect 8392 52640 8444 52649
rect 6920 52572 6972 52624
rect 6184 52436 6236 52488
rect 8208 52479 8260 52488
rect 8208 52445 8217 52479
rect 8217 52445 8251 52479
rect 8251 52445 8260 52479
rect 8208 52436 8260 52445
rect 3010 52198 3062 52250
rect 3074 52198 3126 52250
rect 3138 52198 3190 52250
rect 3202 52198 3254 52250
rect 3266 52198 3318 52250
rect 8010 52198 8062 52250
rect 8074 52198 8126 52250
rect 8138 52198 8190 52250
rect 8202 52198 8254 52250
rect 8266 52198 8318 52250
rect 7932 52096 7984 52148
rect 8116 52096 8168 52148
rect 7932 51960 7984 52012
rect 4436 51935 4488 51944
rect 4436 51901 4445 51935
rect 4445 51901 4479 51935
rect 4479 51901 4488 51935
rect 4436 51892 4488 51901
rect 4712 51935 4764 51944
rect 4712 51901 4721 51935
rect 4721 51901 4755 51935
rect 4755 51901 4764 51935
rect 4712 51892 4764 51901
rect 5724 51756 5776 51808
rect 8392 51799 8444 51808
rect 8392 51765 8401 51799
rect 8401 51765 8435 51799
rect 8435 51765 8444 51799
rect 8392 51756 8444 51765
rect 2350 51654 2402 51706
rect 2414 51654 2466 51706
rect 2478 51654 2530 51706
rect 2542 51654 2594 51706
rect 2606 51654 2658 51706
rect 7350 51654 7402 51706
rect 7414 51654 7466 51706
rect 7478 51654 7530 51706
rect 7542 51654 7594 51706
rect 7606 51654 7658 51706
rect 4712 51552 4764 51604
rect 7104 51552 7156 51604
rect 7380 51552 7432 51604
rect 5724 51459 5776 51468
rect 5724 51425 5733 51459
rect 5733 51425 5767 51459
rect 5767 51425 5776 51459
rect 5724 51416 5776 51425
rect 5908 51459 5960 51468
rect 5908 51425 5917 51459
rect 5917 51425 5951 51459
rect 5951 51425 5960 51459
rect 5908 51416 5960 51425
rect 6736 51459 6788 51468
rect 6736 51425 6745 51459
rect 6745 51425 6779 51459
rect 6779 51425 6788 51459
rect 6736 51416 6788 51425
rect 7012 51416 7064 51468
rect 6184 51348 6236 51400
rect 6460 51391 6512 51400
rect 6460 51357 6469 51391
rect 6469 51357 6503 51391
rect 6503 51357 6512 51391
rect 6460 51348 6512 51357
rect 8116 51348 8168 51400
rect 7932 51212 7984 51264
rect 3010 51110 3062 51162
rect 3074 51110 3126 51162
rect 3138 51110 3190 51162
rect 3202 51110 3254 51162
rect 3266 51110 3318 51162
rect 8010 51110 8062 51162
rect 8074 51110 8126 51162
rect 8138 51110 8190 51162
rect 8202 51110 8254 51162
rect 8266 51110 8318 51162
rect 6460 51008 6512 51060
rect 7932 51008 7984 51060
rect 5724 50915 5776 50924
rect 5724 50881 5733 50915
rect 5733 50881 5767 50915
rect 5767 50881 5776 50915
rect 5724 50872 5776 50881
rect 5816 50847 5868 50856
rect 5816 50813 5825 50847
rect 5825 50813 5859 50847
rect 5859 50813 5868 50847
rect 5816 50804 5868 50813
rect 5908 50847 5960 50856
rect 5908 50813 5917 50847
rect 5917 50813 5951 50847
rect 5951 50813 5960 50847
rect 5908 50804 5960 50813
rect 6920 50804 6972 50856
rect 4896 50668 4948 50720
rect 5724 50668 5776 50720
rect 6552 50668 6604 50720
rect 7104 50668 7156 50720
rect 7380 50668 7432 50720
rect 7840 50668 7892 50720
rect 2350 50566 2402 50618
rect 2414 50566 2466 50618
rect 2478 50566 2530 50618
rect 2542 50566 2594 50618
rect 2606 50566 2658 50618
rect 7350 50566 7402 50618
rect 7414 50566 7466 50618
rect 7478 50566 7530 50618
rect 7542 50566 7594 50618
rect 7606 50566 7658 50618
rect 5816 50464 5868 50516
rect 4896 50328 4948 50380
rect 4436 50260 4488 50312
rect 6460 50303 6512 50312
rect 6460 50269 6469 50303
rect 6469 50269 6503 50303
rect 6503 50269 6512 50303
rect 6460 50260 6512 50269
rect 6552 50260 6604 50312
rect 6736 50303 6788 50312
rect 6736 50269 6745 50303
rect 6745 50269 6779 50303
rect 6779 50269 6788 50303
rect 6736 50260 6788 50269
rect 6920 50124 6972 50176
rect 7932 50124 7984 50176
rect 3010 50022 3062 50074
rect 3074 50022 3126 50074
rect 3138 50022 3190 50074
rect 3202 50022 3254 50074
rect 3266 50022 3318 50074
rect 8010 50022 8062 50074
rect 8074 50022 8126 50074
rect 8138 50022 8190 50074
rect 8202 50022 8254 50074
rect 8266 50022 8318 50074
rect 8392 49963 8444 49972
rect 8392 49929 8401 49963
rect 8401 49929 8435 49963
rect 8435 49929 8444 49963
rect 8392 49920 8444 49929
rect 5540 49784 5592 49836
rect 4436 49716 4488 49768
rect 6552 49716 6604 49768
rect 7012 49648 7064 49700
rect 2350 49478 2402 49530
rect 2414 49478 2466 49530
rect 2478 49478 2530 49530
rect 2542 49478 2594 49530
rect 2606 49478 2658 49530
rect 7350 49478 7402 49530
rect 7414 49478 7466 49530
rect 7478 49478 7530 49530
rect 7542 49478 7594 49530
rect 7606 49478 7658 49530
rect 6460 49376 6512 49428
rect 7472 49376 7524 49428
rect 7932 49376 7984 49428
rect 4436 49172 4488 49224
rect 7104 49240 7156 49292
rect 7012 49215 7064 49224
rect 7012 49181 7021 49215
rect 7021 49181 7055 49215
rect 7055 49181 7064 49215
rect 7012 49172 7064 49181
rect 7748 49172 7800 49224
rect 7932 49172 7984 49224
rect 4988 49147 5040 49156
rect 4988 49113 4997 49147
rect 4997 49113 5031 49147
rect 5031 49113 5040 49147
rect 4988 49104 5040 49113
rect 5908 49036 5960 49088
rect 6644 49036 6696 49088
rect 7288 49036 7340 49088
rect 8392 49079 8444 49088
rect 8392 49045 8401 49079
rect 8401 49045 8435 49079
rect 8435 49045 8444 49079
rect 8392 49036 8444 49045
rect 3010 48934 3062 48986
rect 3074 48934 3126 48986
rect 3138 48934 3190 48986
rect 3202 48934 3254 48986
rect 3266 48934 3318 48986
rect 8010 48934 8062 48986
rect 8074 48934 8126 48986
rect 8138 48934 8190 48986
rect 8202 48934 8254 48986
rect 8266 48934 8318 48986
rect 4988 48832 5040 48884
rect 5816 48875 5868 48884
rect 5816 48841 5825 48875
rect 5825 48841 5859 48875
rect 5859 48841 5868 48875
rect 5816 48832 5868 48841
rect 6644 48832 6696 48884
rect 7288 48832 7340 48884
rect 7472 48764 7524 48816
rect 5908 48671 5960 48680
rect 5908 48637 5917 48671
rect 5917 48637 5951 48671
rect 5951 48637 5960 48671
rect 5908 48628 5960 48637
rect 6000 48671 6052 48680
rect 6000 48637 6009 48671
rect 6009 48637 6043 48671
rect 6043 48637 6052 48671
rect 6000 48628 6052 48637
rect 6552 48628 6604 48680
rect 7104 48628 7156 48680
rect 7656 48628 7708 48680
rect 8024 48492 8076 48544
rect 2350 48390 2402 48442
rect 2414 48390 2466 48442
rect 2478 48390 2530 48442
rect 2542 48390 2594 48442
rect 2606 48390 2658 48442
rect 7350 48390 7402 48442
rect 7414 48390 7466 48442
rect 7478 48390 7530 48442
rect 7542 48390 7594 48442
rect 7606 48390 7658 48442
rect 7748 48288 7800 48340
rect 7104 48220 7156 48272
rect 6000 48195 6052 48204
rect 6000 48161 6009 48195
rect 6009 48161 6043 48195
rect 6043 48161 6052 48195
rect 6000 48152 6052 48161
rect 5908 48084 5960 48136
rect 8024 48084 8076 48136
rect 4896 47948 4948 48000
rect 6184 47948 6236 48000
rect 3010 47846 3062 47898
rect 3074 47846 3126 47898
rect 3138 47846 3190 47898
rect 3202 47846 3254 47898
rect 3266 47846 3318 47898
rect 8010 47846 8062 47898
rect 8074 47846 8126 47898
rect 8138 47846 8190 47898
rect 8202 47846 8254 47898
rect 8266 47846 8318 47898
rect 4896 47744 4948 47796
rect 6092 47676 6144 47728
rect 7104 47676 7156 47728
rect 6460 47651 6512 47660
rect 6460 47617 6469 47651
rect 6469 47617 6503 47651
rect 6503 47617 6512 47651
rect 6460 47608 6512 47617
rect 4436 47583 4488 47592
rect 4436 47549 4445 47583
rect 4445 47549 4479 47583
rect 4479 47549 4488 47583
rect 4436 47540 4488 47549
rect 6552 47540 6604 47592
rect 6184 47447 6236 47456
rect 6184 47413 6193 47447
rect 6193 47413 6227 47447
rect 6227 47413 6236 47447
rect 6184 47404 6236 47413
rect 2350 47302 2402 47354
rect 2414 47302 2466 47354
rect 2478 47302 2530 47354
rect 2542 47302 2594 47354
rect 2606 47302 2658 47354
rect 7350 47302 7402 47354
rect 7414 47302 7466 47354
rect 7478 47302 7530 47354
rect 7542 47302 7594 47354
rect 7606 47302 7658 47354
rect 6460 47200 6512 47252
rect 7012 47200 7064 47252
rect 8392 47243 8444 47252
rect 8392 47209 8401 47243
rect 8401 47209 8435 47243
rect 8435 47209 8444 47243
rect 8392 47200 8444 47209
rect 6000 47107 6052 47116
rect 6000 47073 6009 47107
rect 6009 47073 6043 47107
rect 6043 47073 6052 47107
rect 6000 47064 6052 47073
rect 6184 47064 6236 47116
rect 7380 47107 7432 47116
rect 7380 47073 7389 47107
rect 7389 47073 7423 47107
rect 7423 47073 7432 47107
rect 7380 47064 7432 47073
rect 6460 46996 6512 47048
rect 7104 46996 7156 47048
rect 6092 46928 6144 46980
rect 5448 46903 5500 46912
rect 5448 46869 5457 46903
rect 5457 46869 5491 46903
rect 5491 46869 5500 46903
rect 5448 46860 5500 46869
rect 6184 46860 6236 46912
rect 3010 46758 3062 46810
rect 3074 46758 3126 46810
rect 3138 46758 3190 46810
rect 3202 46758 3254 46810
rect 3266 46758 3318 46810
rect 8010 46758 8062 46810
rect 8074 46758 8126 46810
rect 8138 46758 8190 46810
rect 8202 46758 8254 46810
rect 8266 46758 8318 46810
rect 6460 46588 6512 46640
rect 8024 46588 8076 46640
rect 4436 46495 4488 46504
rect 4436 46461 4445 46495
rect 4445 46461 4479 46495
rect 4479 46461 4488 46495
rect 4436 46452 4488 46461
rect 4712 46495 4764 46504
rect 4712 46461 4721 46495
rect 4721 46461 4755 46495
rect 4755 46461 4764 46495
rect 4712 46452 4764 46461
rect 6184 46495 6236 46504
rect 6184 46461 6193 46495
rect 6193 46461 6227 46495
rect 6227 46461 6236 46495
rect 6184 46452 6236 46461
rect 7380 46495 7432 46504
rect 7380 46461 7389 46495
rect 7389 46461 7423 46495
rect 7423 46461 7432 46495
rect 7380 46452 7432 46461
rect 7840 46452 7892 46504
rect 6828 46359 6880 46368
rect 6828 46325 6837 46359
rect 6837 46325 6871 46359
rect 6871 46325 6880 46359
rect 6828 46316 6880 46325
rect 8392 46359 8444 46368
rect 8392 46325 8401 46359
rect 8401 46325 8435 46359
rect 8435 46325 8444 46359
rect 8392 46316 8444 46325
rect 2350 46214 2402 46266
rect 2414 46214 2466 46266
rect 2478 46214 2530 46266
rect 2542 46214 2594 46266
rect 2606 46214 2658 46266
rect 7350 46214 7402 46266
rect 7414 46214 7466 46266
rect 7478 46214 7530 46266
rect 7542 46214 7594 46266
rect 7606 46214 7658 46266
rect 4712 46112 4764 46164
rect 6828 46112 6880 46164
rect 6000 45976 6052 46028
rect 5448 45908 5500 45960
rect 6184 45908 6236 45960
rect 6552 45908 6604 45960
rect 8024 45908 8076 45960
rect 5632 45772 5684 45824
rect 5724 45772 5776 45824
rect 6092 45772 6144 45824
rect 3010 45670 3062 45722
rect 3074 45670 3126 45722
rect 3138 45670 3190 45722
rect 3202 45670 3254 45722
rect 3266 45670 3318 45722
rect 8010 45670 8062 45722
rect 8074 45670 8126 45722
rect 8138 45670 8190 45722
rect 8202 45670 8254 45722
rect 8266 45670 8318 45722
rect 6092 45611 6144 45620
rect 6092 45577 6101 45611
rect 6101 45577 6135 45611
rect 6135 45577 6144 45611
rect 6092 45568 6144 45577
rect 6460 45432 6512 45484
rect 6920 45432 6972 45484
rect 7104 45432 7156 45484
rect 4620 45407 4672 45416
rect 4620 45373 4629 45407
rect 4629 45373 4663 45407
rect 4663 45373 4672 45407
rect 4620 45364 4672 45373
rect 7840 45364 7892 45416
rect 4436 45228 4488 45280
rect 6920 45271 6972 45280
rect 6920 45237 6929 45271
rect 6929 45237 6963 45271
rect 6963 45237 6972 45271
rect 6920 45228 6972 45237
rect 2350 45126 2402 45178
rect 2414 45126 2466 45178
rect 2478 45126 2530 45178
rect 2542 45126 2594 45178
rect 2606 45126 2658 45178
rect 7350 45126 7402 45178
rect 7414 45126 7466 45178
rect 7478 45126 7530 45178
rect 7542 45126 7594 45178
rect 7606 45126 7658 45178
rect 4620 45024 4672 45076
rect 5632 44820 5684 44872
rect 6552 44820 6604 44872
rect 8024 44820 8076 44872
rect 7196 44684 7248 44736
rect 3010 44582 3062 44634
rect 3074 44582 3126 44634
rect 3138 44582 3190 44634
rect 3202 44582 3254 44634
rect 3266 44582 3318 44634
rect 8010 44582 8062 44634
rect 8074 44582 8126 44634
rect 8138 44582 8190 44634
rect 8202 44582 8254 44634
rect 8266 44582 8318 44634
rect 6920 44480 6972 44532
rect 7196 44480 7248 44532
rect 8392 44523 8444 44532
rect 8392 44489 8401 44523
rect 8401 44489 8435 44523
rect 8435 44489 8444 44523
rect 8392 44480 8444 44489
rect 5356 44387 5408 44396
rect 5356 44353 5365 44387
rect 5365 44353 5399 44387
rect 5399 44353 5408 44387
rect 5356 44344 5408 44353
rect 5172 44183 5224 44192
rect 5172 44149 5181 44183
rect 5181 44149 5215 44183
rect 5215 44149 5224 44183
rect 5172 44140 5224 44149
rect 2350 44038 2402 44090
rect 2414 44038 2466 44090
rect 2478 44038 2530 44090
rect 2542 44038 2594 44090
rect 2606 44038 2658 44090
rect 7350 44038 7402 44090
rect 7414 44038 7466 44090
rect 7478 44038 7530 44090
rect 7542 44038 7594 44090
rect 7606 44038 7658 44090
rect 6276 43936 6328 43988
rect 5172 43843 5224 43852
rect 5172 43809 5181 43843
rect 5181 43809 5215 43843
rect 5215 43809 5224 43843
rect 5172 43800 5224 43809
rect 4436 43732 4488 43784
rect 6460 43732 6512 43784
rect 7932 43596 7984 43648
rect 8852 43596 8904 43648
rect 3010 43494 3062 43546
rect 3074 43494 3126 43546
rect 3138 43494 3190 43546
rect 3202 43494 3254 43546
rect 3266 43494 3318 43546
rect 8010 43494 8062 43546
rect 8074 43494 8126 43546
rect 8138 43494 8190 43546
rect 8202 43494 8254 43546
rect 8266 43494 8318 43546
rect 5356 43435 5408 43444
rect 5356 43401 5365 43435
rect 5365 43401 5399 43435
rect 5399 43401 5408 43435
rect 5356 43392 5408 43401
rect 6276 43392 6328 43444
rect 6920 43392 6972 43444
rect 7104 43392 7156 43444
rect 6184 43256 6236 43308
rect 7104 43256 7156 43308
rect 7196 43256 7248 43308
rect 6000 43231 6052 43240
rect 6000 43197 6009 43231
rect 6009 43197 6043 43231
rect 6043 43197 6052 43231
rect 6000 43188 6052 43197
rect 6920 43052 6972 43104
rect 2350 42950 2402 43002
rect 2414 42950 2466 43002
rect 2478 42950 2530 43002
rect 2542 42950 2594 43002
rect 2606 42950 2658 43002
rect 7350 42950 7402 43002
rect 7414 42950 7466 43002
rect 7478 42950 7530 43002
rect 7542 42950 7594 43002
rect 7606 42950 7658 43002
rect 6920 42848 6972 42900
rect 6552 42755 6604 42764
rect 6552 42721 6561 42755
rect 6561 42721 6595 42755
rect 6595 42721 6604 42755
rect 6552 42712 6604 42721
rect 4436 42644 4488 42696
rect 6460 42644 6512 42696
rect 4988 42619 5040 42628
rect 4988 42585 4997 42619
rect 4997 42585 5031 42619
rect 5031 42585 5040 42619
rect 4988 42576 5040 42585
rect 6828 42576 6880 42628
rect 7104 42508 7156 42560
rect 7840 42508 7892 42560
rect 3010 42406 3062 42458
rect 3074 42406 3126 42458
rect 3138 42406 3190 42458
rect 3202 42406 3254 42458
rect 3266 42406 3318 42458
rect 8010 42406 8062 42458
rect 8074 42406 8126 42458
rect 8138 42406 8190 42458
rect 8202 42406 8254 42458
rect 8266 42406 8318 42458
rect 4988 42304 5040 42356
rect 5908 42236 5960 42288
rect 7104 42304 7156 42356
rect 7196 42304 7248 42356
rect 6184 42236 6236 42288
rect 7840 42236 7892 42288
rect 7932 42236 7984 42288
rect 6920 42100 6972 42152
rect 8392 42032 8444 42084
rect 2350 41862 2402 41914
rect 2414 41862 2466 41914
rect 2478 41862 2530 41914
rect 2542 41862 2594 41914
rect 2606 41862 2658 41914
rect 7350 41862 7402 41914
rect 7414 41862 7466 41914
rect 7478 41862 7530 41914
rect 7542 41862 7594 41914
rect 7606 41862 7658 41914
rect 5908 41760 5960 41812
rect 6736 41556 6788 41608
rect 6920 41556 6972 41608
rect 6184 41531 6236 41540
rect 6184 41497 6193 41531
rect 6193 41497 6227 41531
rect 6227 41497 6236 41531
rect 6184 41488 6236 41497
rect 7840 41488 7892 41540
rect 7748 41420 7800 41472
rect 3010 41318 3062 41370
rect 3074 41318 3126 41370
rect 3138 41318 3190 41370
rect 3202 41318 3254 41370
rect 3266 41318 3318 41370
rect 8010 41318 8062 41370
rect 8074 41318 8126 41370
rect 8138 41318 8190 41370
rect 8202 41318 8254 41370
rect 8266 41318 8318 41370
rect 6092 41216 6144 41268
rect 6920 41148 6972 41200
rect 7104 41148 7156 41200
rect 4436 41123 4488 41132
rect 4436 41089 4445 41123
rect 4445 41089 4479 41123
rect 4479 41089 4488 41123
rect 4436 41080 4488 41089
rect 6460 41123 6512 41132
rect 6460 41089 6469 41123
rect 6469 41089 6503 41123
rect 6503 41089 6512 41123
rect 6460 41080 6512 41089
rect 4712 41055 4764 41064
rect 4712 41021 4721 41055
rect 4721 41021 4755 41055
rect 4755 41021 4764 41055
rect 4712 41012 4764 41021
rect 6920 40876 6972 40928
rect 8392 40919 8444 40928
rect 8392 40885 8401 40919
rect 8401 40885 8435 40919
rect 8435 40885 8444 40919
rect 8392 40876 8444 40885
rect 2350 40774 2402 40826
rect 2414 40774 2466 40826
rect 2478 40774 2530 40826
rect 2542 40774 2594 40826
rect 2606 40774 2658 40826
rect 7350 40774 7402 40826
rect 7414 40774 7466 40826
rect 7478 40774 7530 40826
rect 7542 40774 7594 40826
rect 7606 40774 7658 40826
rect 4712 40672 4764 40724
rect 4804 40511 4856 40520
rect 4804 40477 4813 40511
rect 4813 40477 4847 40511
rect 4847 40477 4856 40511
rect 4804 40468 4856 40477
rect 7012 40536 7064 40588
rect 6736 40511 6788 40520
rect 6736 40477 6745 40511
rect 6745 40477 6779 40511
rect 6779 40477 6788 40511
rect 6736 40468 6788 40477
rect 6920 40400 6972 40452
rect 7104 40400 7156 40452
rect 5540 40332 5592 40384
rect 6828 40332 6880 40384
rect 3010 40230 3062 40282
rect 3074 40230 3126 40282
rect 3138 40230 3190 40282
rect 3202 40230 3254 40282
rect 3266 40230 3318 40282
rect 8010 40230 8062 40282
rect 8074 40230 8126 40282
rect 8138 40230 8190 40282
rect 8202 40230 8254 40282
rect 8266 40230 8318 40282
rect 4804 40128 4856 40180
rect 6092 40128 6144 40180
rect 6368 40128 6420 40180
rect 6460 40128 6512 40180
rect 5632 40103 5684 40112
rect 5632 40069 5641 40103
rect 5641 40069 5675 40103
rect 5675 40069 5684 40103
rect 5632 40060 5684 40069
rect 5908 39967 5960 39976
rect 5908 39933 5917 39967
rect 5917 39933 5951 39967
rect 5951 39933 5960 39967
rect 5908 39924 5960 39933
rect 6276 39924 6328 39976
rect 7748 39924 7800 39976
rect 6552 39831 6604 39840
rect 6552 39797 6561 39831
rect 6561 39797 6595 39831
rect 6595 39797 6604 39831
rect 6552 39788 6604 39797
rect 2350 39686 2402 39738
rect 2414 39686 2466 39738
rect 2478 39686 2530 39738
rect 2542 39686 2594 39738
rect 2606 39686 2658 39738
rect 7350 39686 7402 39738
rect 7414 39686 7466 39738
rect 7478 39686 7530 39738
rect 7542 39686 7594 39738
rect 7606 39686 7658 39738
rect 4436 39380 4488 39432
rect 6736 39423 6788 39432
rect 6736 39389 6745 39423
rect 6745 39389 6779 39423
rect 6779 39389 6788 39423
rect 6736 39380 6788 39389
rect 4988 39355 5040 39364
rect 4988 39321 4997 39355
rect 4997 39321 5031 39355
rect 5031 39321 5040 39355
rect 4988 39312 5040 39321
rect 6552 39312 6604 39364
rect 5908 39244 5960 39296
rect 7104 39312 7156 39364
rect 7656 39244 7708 39296
rect 3010 39142 3062 39194
rect 3074 39142 3126 39194
rect 3138 39142 3190 39194
rect 3202 39142 3254 39194
rect 3266 39142 3318 39194
rect 8010 39142 8062 39194
rect 8074 39142 8126 39194
rect 8138 39142 8190 39194
rect 8202 39142 8254 39194
rect 8266 39142 8318 39194
rect 4988 39040 5040 39092
rect 6276 38972 6328 39024
rect 5908 38947 5960 38956
rect 5908 38913 5917 38947
rect 5917 38913 5951 38947
rect 5951 38913 5960 38947
rect 5908 38904 5960 38913
rect 7656 39040 7708 39092
rect 8392 39083 8444 39092
rect 8392 39049 8401 39083
rect 8401 39049 8435 39083
rect 8435 39049 8444 39083
rect 8392 39040 8444 39049
rect 6092 38879 6144 38888
rect 6092 38845 6101 38879
rect 6101 38845 6135 38879
rect 6135 38845 6144 38879
rect 6092 38836 6144 38845
rect 7196 38768 7248 38820
rect 7748 38768 7800 38820
rect 2350 38598 2402 38650
rect 2414 38598 2466 38650
rect 2478 38598 2530 38650
rect 2542 38598 2594 38650
rect 2606 38598 2658 38650
rect 7350 38598 7402 38650
rect 7414 38598 7466 38650
rect 7478 38598 7530 38650
rect 7542 38598 7594 38650
rect 7606 38598 7658 38650
rect 7104 38360 7156 38412
rect 4436 38292 4488 38344
rect 6000 38292 6052 38344
rect 7748 38292 7800 38344
rect 4896 38267 4948 38276
rect 4896 38233 4905 38267
rect 4905 38233 4939 38267
rect 4939 38233 4948 38267
rect 4896 38224 4948 38233
rect 6552 38267 6604 38276
rect 6552 38233 6561 38267
rect 6561 38233 6595 38267
rect 6595 38233 6604 38267
rect 6552 38224 6604 38233
rect 5816 38156 5868 38208
rect 8392 38199 8444 38208
rect 8392 38165 8401 38199
rect 8401 38165 8435 38199
rect 8435 38165 8444 38199
rect 8392 38156 8444 38165
rect 3010 38054 3062 38106
rect 3074 38054 3126 38106
rect 3138 38054 3190 38106
rect 3202 38054 3254 38106
rect 3266 38054 3318 38106
rect 8010 38054 8062 38106
rect 8074 38054 8126 38106
rect 8138 38054 8190 38106
rect 8202 38054 8254 38106
rect 8266 38054 8318 38106
rect 4896 37952 4948 38004
rect 5908 37952 5960 38004
rect 8024 37884 8076 37936
rect 6460 37859 6512 37868
rect 6460 37825 6469 37859
rect 6469 37825 6503 37859
rect 6503 37825 6512 37859
rect 6460 37816 6512 37825
rect 5908 37791 5960 37800
rect 5908 37757 5917 37791
rect 5917 37757 5951 37791
rect 5951 37757 5960 37791
rect 5908 37748 5960 37757
rect 6092 37791 6144 37800
rect 6092 37757 6101 37791
rect 6101 37757 6135 37791
rect 6135 37757 6144 37791
rect 6092 37748 6144 37757
rect 6736 37791 6788 37800
rect 6736 37757 6745 37791
rect 6745 37757 6779 37791
rect 6779 37757 6788 37791
rect 6736 37748 6788 37757
rect 7104 37612 7156 37664
rect 7748 37612 7800 37664
rect 2350 37510 2402 37562
rect 2414 37510 2466 37562
rect 2478 37510 2530 37562
rect 2542 37510 2594 37562
rect 2606 37510 2658 37562
rect 7350 37510 7402 37562
rect 7414 37510 7466 37562
rect 7478 37510 7530 37562
rect 7542 37510 7594 37562
rect 7606 37510 7658 37562
rect 6460 37408 6512 37460
rect 6092 37272 6144 37324
rect 7196 37272 7248 37324
rect 5080 37111 5132 37120
rect 5080 37077 5089 37111
rect 5089 37077 5123 37111
rect 5123 37077 5132 37111
rect 5080 37068 5132 37077
rect 7104 37247 7156 37256
rect 7104 37213 7113 37247
rect 7113 37213 7147 37247
rect 7147 37213 7156 37247
rect 7104 37204 7156 37213
rect 5908 37136 5960 37188
rect 6184 37068 6236 37120
rect 3010 36966 3062 37018
rect 3074 36966 3126 37018
rect 3138 36966 3190 37018
rect 3202 36966 3254 37018
rect 3266 36966 3318 37018
rect 8010 36966 8062 37018
rect 8074 36966 8126 37018
rect 8138 36966 8190 37018
rect 8202 36966 8254 37018
rect 8266 36966 8318 37018
rect 5080 36864 5132 36916
rect 6184 36907 6236 36916
rect 6184 36873 6193 36907
rect 6193 36873 6227 36907
rect 6227 36873 6236 36907
rect 6184 36864 6236 36873
rect 7932 36864 7984 36916
rect 4436 36703 4488 36712
rect 4436 36669 4445 36703
rect 4445 36669 4479 36703
rect 4479 36669 4488 36703
rect 4436 36660 4488 36669
rect 6460 36771 6512 36780
rect 6460 36737 6469 36771
rect 6469 36737 6503 36771
rect 6503 36737 6512 36771
rect 6460 36728 6512 36737
rect 6736 36703 6788 36712
rect 6736 36669 6745 36703
rect 6745 36669 6779 36703
rect 6779 36669 6788 36703
rect 6736 36660 6788 36669
rect 6000 36592 6052 36644
rect 7748 36660 7800 36712
rect 2350 36422 2402 36474
rect 2414 36422 2466 36474
rect 2478 36422 2530 36474
rect 2542 36422 2594 36474
rect 2606 36422 2658 36474
rect 7350 36422 7402 36474
rect 7414 36422 7466 36474
rect 7478 36422 7530 36474
rect 7542 36422 7594 36474
rect 7606 36422 7658 36474
rect 6460 36320 6512 36372
rect 8392 36363 8444 36372
rect 8392 36329 8401 36363
rect 8401 36329 8435 36363
rect 8435 36329 8444 36363
rect 8392 36320 8444 36329
rect 6184 36184 6236 36236
rect 7196 36227 7248 36236
rect 7196 36193 7205 36227
rect 7205 36193 7239 36227
rect 7239 36193 7248 36227
rect 7196 36184 7248 36193
rect 3010 35878 3062 35930
rect 3074 35878 3126 35930
rect 3138 35878 3190 35930
rect 3202 35878 3254 35930
rect 3266 35878 3318 35930
rect 8010 35878 8062 35930
rect 8074 35878 8126 35930
rect 8138 35878 8190 35930
rect 8202 35878 8254 35930
rect 8266 35878 8318 35930
rect 6184 35776 6236 35828
rect 8024 35640 8076 35692
rect 5908 35615 5960 35624
rect 5908 35581 5917 35615
rect 5917 35581 5951 35615
rect 5951 35581 5960 35615
rect 5908 35572 5960 35581
rect 6092 35615 6144 35624
rect 6092 35581 6101 35615
rect 6101 35581 6135 35615
rect 6135 35581 6144 35615
rect 6092 35572 6144 35581
rect 4988 35436 5040 35488
rect 8392 35479 8444 35488
rect 8392 35445 8401 35479
rect 8401 35445 8435 35479
rect 8435 35445 8444 35479
rect 8392 35436 8444 35445
rect 2350 35334 2402 35386
rect 2414 35334 2466 35386
rect 2478 35334 2530 35386
rect 2542 35334 2594 35386
rect 2606 35334 2658 35386
rect 7350 35334 7402 35386
rect 7414 35334 7466 35386
rect 7478 35334 7530 35386
rect 7542 35334 7594 35386
rect 7606 35334 7658 35386
rect 5908 35232 5960 35284
rect 4988 35096 5040 35148
rect 4436 35028 4488 35080
rect 6460 35071 6512 35080
rect 6460 35037 6469 35071
rect 6469 35037 6503 35071
rect 6503 35037 6512 35071
rect 6460 35028 6512 35037
rect 6736 35071 6788 35080
rect 6736 35037 6745 35071
rect 6745 35037 6779 35071
rect 6779 35037 6788 35071
rect 6736 35028 6788 35037
rect 6184 34960 6236 35012
rect 4804 34892 4856 34944
rect 7288 34960 7340 35012
rect 7104 34892 7156 34944
rect 8024 34892 8076 34944
rect 3010 34790 3062 34842
rect 3074 34790 3126 34842
rect 3138 34790 3190 34842
rect 3202 34790 3254 34842
rect 3266 34790 3318 34842
rect 8010 34790 8062 34842
rect 8074 34790 8126 34842
rect 8138 34790 8190 34842
rect 8202 34790 8254 34842
rect 8266 34790 8318 34842
rect 5448 34552 5500 34604
rect 6828 34595 6880 34604
rect 6828 34561 6837 34595
rect 6837 34561 6871 34595
rect 6871 34561 6880 34595
rect 6828 34552 6880 34561
rect 4804 34484 4856 34536
rect 6736 34484 6788 34536
rect 5632 34391 5684 34400
rect 5632 34357 5641 34391
rect 5641 34357 5675 34391
rect 5675 34357 5684 34391
rect 5632 34348 5684 34357
rect 2350 34246 2402 34298
rect 2414 34246 2466 34298
rect 2478 34246 2530 34298
rect 2542 34246 2594 34298
rect 2606 34246 2658 34298
rect 7350 34246 7402 34298
rect 7414 34246 7466 34298
rect 7478 34246 7530 34298
rect 7542 34246 7594 34298
rect 7606 34246 7658 34298
rect 5632 34144 5684 34196
rect 4804 34076 4856 34128
rect 7012 34008 7064 34060
rect 7380 34008 7432 34060
rect 6184 33940 6236 33992
rect 6552 33847 6604 33856
rect 6552 33813 6561 33847
rect 6561 33813 6595 33847
rect 6595 33813 6604 33847
rect 6552 33804 6604 33813
rect 6736 33804 6788 33856
rect 7012 33915 7064 33924
rect 7012 33881 7021 33915
rect 7021 33881 7055 33915
rect 7055 33881 7064 33915
rect 7012 33872 7064 33881
rect 7196 33804 7248 33856
rect 7932 33804 7984 33856
rect 3010 33702 3062 33754
rect 3074 33702 3126 33754
rect 3138 33702 3190 33754
rect 3202 33702 3254 33754
rect 3266 33702 3318 33754
rect 8010 33702 8062 33754
rect 8074 33702 8126 33754
rect 8138 33702 8190 33754
rect 8202 33702 8254 33754
rect 8266 33702 8318 33754
rect 5448 33643 5500 33652
rect 5448 33609 5457 33643
rect 5457 33609 5491 33643
rect 5491 33609 5500 33643
rect 5448 33600 5500 33609
rect 5816 33643 5868 33652
rect 5816 33609 5825 33643
rect 5825 33609 5859 33643
rect 5859 33609 5868 33643
rect 5816 33600 5868 33609
rect 6460 33600 6512 33652
rect 7104 33643 7156 33652
rect 7104 33609 7113 33643
rect 7113 33609 7147 33643
rect 7147 33609 7156 33643
rect 7104 33600 7156 33609
rect 7932 33643 7984 33652
rect 7932 33609 7941 33643
rect 7941 33609 7975 33643
rect 7975 33609 7984 33643
rect 7932 33600 7984 33609
rect 6552 33532 6604 33584
rect 6092 33439 6144 33448
rect 6092 33405 6101 33439
rect 6101 33405 6135 33439
rect 6135 33405 6144 33439
rect 6092 33396 6144 33405
rect 7380 33439 7432 33448
rect 7380 33405 7389 33439
rect 7389 33405 7423 33439
rect 7423 33405 7432 33439
rect 7380 33396 7432 33405
rect 8024 33396 8076 33448
rect 7196 33260 7248 33312
rect 2350 33158 2402 33210
rect 2414 33158 2466 33210
rect 2478 33158 2530 33210
rect 2542 33158 2594 33210
rect 2606 33158 2658 33210
rect 7350 33158 7402 33210
rect 7414 33158 7466 33210
rect 7478 33158 7530 33210
rect 7542 33158 7594 33210
rect 7606 33158 7658 33210
rect 7012 33099 7064 33108
rect 7012 33065 7021 33099
rect 7021 33065 7055 33099
rect 7055 33065 7064 33099
rect 7012 33056 7064 33065
rect 7748 33056 7800 33108
rect 7932 33056 7984 33108
rect 7196 32895 7248 32904
rect 7196 32861 7205 32895
rect 7205 32861 7239 32895
rect 7239 32861 7248 32895
rect 7196 32852 7248 32861
rect 7748 32784 7800 32836
rect 8668 32716 8720 32768
rect 3010 32614 3062 32666
rect 3074 32614 3126 32666
rect 3138 32614 3190 32666
rect 3202 32614 3254 32666
rect 3266 32614 3318 32666
rect 8010 32614 8062 32666
rect 8074 32614 8126 32666
rect 8138 32614 8190 32666
rect 8202 32614 8254 32666
rect 8266 32614 8318 32666
rect 7104 32444 7156 32496
rect 6460 32419 6512 32428
rect 6460 32385 6469 32419
rect 6469 32385 6503 32419
rect 6503 32385 6512 32419
rect 6460 32376 6512 32385
rect 6552 32376 6604 32428
rect 4712 32351 4764 32360
rect 4712 32317 4721 32351
rect 4721 32317 4755 32351
rect 4755 32317 4764 32351
rect 4712 32308 4764 32317
rect 6736 32351 6788 32360
rect 6736 32317 6745 32351
rect 6745 32317 6779 32351
rect 6779 32317 6788 32351
rect 6736 32308 6788 32317
rect 4804 32172 4856 32224
rect 6184 32215 6236 32224
rect 6184 32181 6193 32215
rect 6193 32181 6227 32215
rect 6227 32181 6236 32215
rect 6184 32172 6236 32181
rect 7104 32172 7156 32224
rect 7748 32172 7800 32224
rect 2350 32070 2402 32122
rect 2414 32070 2466 32122
rect 2478 32070 2530 32122
rect 2542 32070 2594 32122
rect 2606 32070 2658 32122
rect 7350 32070 7402 32122
rect 7414 32070 7466 32122
rect 7478 32070 7530 32122
rect 7542 32070 7594 32122
rect 7606 32070 7658 32122
rect 4712 31968 4764 32020
rect 6460 31968 6512 32020
rect 6000 31832 6052 31884
rect 7748 31832 7800 31884
rect 7932 31832 7984 31884
rect 6920 31764 6972 31816
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 6184 31628 6236 31680
rect 3010 31526 3062 31578
rect 3074 31526 3126 31578
rect 3138 31526 3190 31578
rect 3202 31526 3254 31578
rect 3266 31526 3318 31578
rect 8010 31526 8062 31578
rect 8074 31526 8126 31578
rect 8138 31526 8190 31578
rect 8202 31526 8254 31578
rect 8266 31526 8318 31578
rect 8024 31356 8076 31408
rect 6460 31331 6512 31340
rect 6460 31297 6469 31331
rect 6469 31297 6503 31331
rect 6503 31297 6512 31331
rect 6460 31288 6512 31297
rect 6736 31263 6788 31272
rect 6736 31229 6745 31263
rect 6745 31229 6779 31263
rect 6779 31229 6788 31263
rect 6736 31220 6788 31229
rect 2350 30982 2402 31034
rect 2414 30982 2466 31034
rect 2478 30982 2530 31034
rect 2542 30982 2594 31034
rect 2606 30982 2658 31034
rect 7350 30982 7402 31034
rect 7414 30982 7466 31034
rect 7478 30982 7530 31034
rect 7542 30982 7594 31034
rect 7606 30982 7658 31034
rect 6460 30880 6512 30932
rect 8024 30880 8076 30932
rect 8392 30923 8444 30932
rect 8392 30889 8401 30923
rect 8401 30889 8435 30923
rect 8435 30889 8444 30923
rect 8392 30880 8444 30889
rect 4804 30787 4856 30796
rect 4804 30753 4813 30787
rect 4813 30753 4847 30787
rect 4847 30753 4856 30787
rect 4804 30744 4856 30753
rect 6460 30744 6512 30796
rect 7748 30744 7800 30796
rect 6552 30676 6604 30728
rect 5080 30651 5132 30660
rect 5080 30617 5089 30651
rect 5089 30617 5123 30651
rect 5123 30617 5132 30651
rect 5080 30608 5132 30617
rect 6644 30540 6696 30592
rect 3010 30438 3062 30490
rect 3074 30438 3126 30490
rect 3138 30438 3190 30490
rect 3202 30438 3254 30490
rect 3266 30438 3318 30490
rect 8010 30438 8062 30490
rect 8074 30438 8126 30490
rect 8138 30438 8190 30490
rect 8202 30438 8254 30490
rect 8266 30438 8318 30490
rect 5080 30336 5132 30388
rect 6184 30336 6236 30388
rect 6460 30336 6512 30388
rect 6092 30268 6144 30320
rect 6644 30132 6696 30184
rect 8392 30039 8444 30048
rect 8392 30005 8401 30039
rect 8401 30005 8435 30039
rect 8435 30005 8444 30039
rect 8392 29996 8444 30005
rect 2350 29894 2402 29946
rect 2414 29894 2466 29946
rect 2478 29894 2530 29946
rect 2542 29894 2594 29946
rect 2606 29894 2658 29946
rect 7350 29894 7402 29946
rect 7414 29894 7466 29946
rect 7478 29894 7530 29946
rect 7542 29894 7594 29946
rect 7606 29894 7658 29946
rect 6092 29699 6144 29708
rect 6092 29665 6101 29699
rect 6101 29665 6135 29699
rect 6135 29665 6144 29699
rect 6092 29656 6144 29665
rect 6276 29656 6328 29708
rect 6460 29631 6512 29640
rect 6460 29597 6469 29631
rect 6469 29597 6503 29631
rect 6503 29597 6512 29631
rect 6460 29588 6512 29597
rect 6736 29631 6788 29640
rect 6736 29597 6745 29631
rect 6745 29597 6779 29631
rect 6779 29597 6788 29631
rect 6736 29588 6788 29597
rect 8024 29588 8076 29640
rect 5264 29452 5316 29504
rect 5908 29495 5960 29504
rect 5908 29461 5917 29495
rect 5917 29461 5951 29495
rect 5951 29461 5960 29495
rect 5908 29452 5960 29461
rect 3010 29350 3062 29402
rect 3074 29350 3126 29402
rect 3138 29350 3190 29402
rect 3202 29350 3254 29402
rect 3266 29350 3318 29402
rect 8010 29350 8062 29402
rect 8074 29350 8126 29402
rect 8138 29350 8190 29402
rect 8202 29350 8254 29402
rect 8266 29350 8318 29402
rect 5264 29248 5316 29300
rect 6460 29248 6512 29300
rect 6644 29180 6696 29232
rect 5908 29155 5960 29164
rect 5908 29121 5917 29155
rect 5917 29121 5951 29155
rect 5951 29121 5960 29155
rect 5908 29112 5960 29121
rect 6092 29087 6144 29096
rect 6092 29053 6101 29087
rect 6101 29053 6135 29087
rect 6135 29053 6144 29087
rect 6092 29044 6144 29053
rect 6552 29044 6604 29096
rect 7196 28976 7248 29028
rect 7748 29044 7800 29096
rect 4712 28908 4764 28960
rect 5172 28951 5224 28960
rect 5172 28917 5181 28951
rect 5181 28917 5215 28951
rect 5215 28917 5224 28951
rect 5172 28908 5224 28917
rect 2350 28806 2402 28858
rect 2414 28806 2466 28858
rect 2478 28806 2530 28858
rect 2542 28806 2594 28858
rect 2606 28806 2658 28858
rect 7350 28806 7402 28858
rect 7414 28806 7466 28858
rect 7478 28806 7530 28858
rect 7542 28806 7594 28858
rect 7606 28806 7658 28858
rect 4804 28611 4856 28620
rect 4804 28577 4813 28611
rect 4813 28577 4847 28611
rect 4847 28577 4856 28611
rect 4804 28568 4856 28577
rect 5172 28568 5224 28620
rect 6092 28500 6144 28552
rect 7104 28568 7156 28620
rect 6736 28543 6788 28552
rect 6736 28509 6745 28543
rect 6745 28509 6779 28543
rect 6779 28509 6788 28543
rect 6736 28500 6788 28509
rect 8024 28500 8076 28552
rect 7012 28475 7064 28484
rect 7012 28441 7021 28475
rect 7021 28441 7055 28475
rect 7055 28441 7064 28475
rect 7012 28432 7064 28441
rect 6552 28407 6604 28416
rect 6552 28373 6561 28407
rect 6561 28373 6595 28407
rect 6595 28373 6604 28407
rect 6552 28364 6604 28373
rect 3010 28262 3062 28314
rect 3074 28262 3126 28314
rect 3138 28262 3190 28314
rect 3202 28262 3254 28314
rect 3266 28262 3318 28314
rect 8010 28262 8062 28314
rect 8074 28262 8126 28314
rect 8138 28262 8190 28314
rect 8202 28262 8254 28314
rect 8266 28262 8318 28314
rect 4804 28160 4856 28212
rect 6092 28160 6144 28212
rect 6276 28160 6328 28212
rect 7012 28160 7064 28212
rect 8392 28203 8444 28212
rect 8392 28169 8401 28203
rect 8401 28169 8435 28203
rect 8435 28169 8444 28203
rect 8392 28160 8444 28169
rect 6552 28092 6604 28144
rect 4436 28067 4488 28076
rect 4436 28033 4445 28067
rect 4445 28033 4479 28067
rect 4479 28033 4488 28067
rect 4436 28024 4488 28033
rect 4712 27999 4764 28008
rect 4712 27965 4721 27999
rect 4721 27965 4755 27999
rect 4755 27965 4764 27999
rect 4712 27956 4764 27965
rect 7196 27956 7248 28008
rect 2350 27718 2402 27770
rect 2414 27718 2466 27770
rect 2478 27718 2530 27770
rect 2542 27718 2594 27770
rect 2606 27718 2658 27770
rect 7350 27718 7402 27770
rect 7414 27718 7466 27770
rect 7478 27718 7530 27770
rect 7542 27718 7594 27770
rect 7606 27718 7658 27770
rect 7932 27344 7984 27396
rect 7840 27276 7892 27328
rect 8392 27276 8444 27328
rect 8852 27276 8904 27328
rect 3010 27174 3062 27226
rect 3074 27174 3126 27226
rect 3138 27174 3190 27226
rect 3202 27174 3254 27226
rect 3266 27174 3318 27226
rect 8010 27174 8062 27226
rect 8074 27174 8126 27226
rect 8138 27174 8190 27226
rect 8202 27174 8254 27226
rect 8266 27174 8318 27226
rect 8392 27072 8444 27124
rect 7196 26936 7248 26988
rect 5724 26868 5776 26920
rect 6184 26868 6236 26920
rect 6920 26911 6972 26920
rect 6920 26877 6929 26911
rect 6929 26877 6963 26911
rect 6963 26877 6972 26911
rect 6920 26868 6972 26877
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 6368 26775 6420 26784
rect 6368 26741 6377 26775
rect 6377 26741 6411 26775
rect 6411 26741 6420 26775
rect 6368 26732 6420 26741
rect 7932 26732 7984 26784
rect 2350 26630 2402 26682
rect 2414 26630 2466 26682
rect 2478 26630 2530 26682
rect 2542 26630 2594 26682
rect 2606 26630 2658 26682
rect 7350 26630 7402 26682
rect 7414 26630 7466 26682
rect 7478 26630 7530 26682
rect 7542 26630 7594 26682
rect 7606 26630 7658 26682
rect 5724 26528 5776 26580
rect 6920 26528 6972 26580
rect 7748 26571 7800 26580
rect 7748 26537 7757 26571
rect 7757 26537 7791 26571
rect 7791 26537 7800 26571
rect 7748 26528 7800 26537
rect 4436 26392 4488 26444
rect 6736 26392 6788 26444
rect 6920 26392 6972 26444
rect 6184 26299 6236 26308
rect 6184 26265 6193 26299
rect 6193 26265 6227 26299
rect 6227 26265 6236 26299
rect 6184 26256 6236 26265
rect 7748 26324 7800 26376
rect 8024 26324 8076 26376
rect 3010 26086 3062 26138
rect 3074 26086 3126 26138
rect 3138 26086 3190 26138
rect 3202 26086 3254 26138
rect 3266 26086 3318 26138
rect 8010 26086 8062 26138
rect 8074 26086 8126 26138
rect 8138 26086 8190 26138
rect 8202 26086 8254 26138
rect 8266 26086 8318 26138
rect 6092 25984 6144 26036
rect 6184 25984 6236 26036
rect 7932 25984 7984 26036
rect 7012 25848 7064 25900
rect 6368 25712 6420 25764
rect 6644 25687 6696 25696
rect 6644 25653 6653 25687
rect 6653 25653 6687 25687
rect 6687 25653 6696 25687
rect 6644 25644 6696 25653
rect 6736 25644 6788 25696
rect 2350 25542 2402 25594
rect 2414 25542 2466 25594
rect 2478 25542 2530 25594
rect 2542 25542 2594 25594
rect 2606 25542 2658 25594
rect 7350 25542 7402 25594
rect 7414 25542 7466 25594
rect 7478 25542 7530 25594
rect 7542 25542 7594 25594
rect 7606 25542 7658 25594
rect 6644 25440 6696 25492
rect 7196 25440 7248 25492
rect 7840 25304 7892 25356
rect 6644 25100 6696 25152
rect 3010 24998 3062 25050
rect 3074 24998 3126 25050
rect 3138 24998 3190 25050
rect 3202 24998 3254 25050
rect 3266 24998 3318 25050
rect 8010 24998 8062 25050
rect 8074 24998 8126 25050
rect 8138 24998 8190 25050
rect 8202 24998 8254 25050
rect 8266 24998 8318 25050
rect 6736 24896 6788 24948
rect 7012 24896 7064 24948
rect 6644 24556 6696 24608
rect 8392 24556 8444 24608
rect 2350 24454 2402 24506
rect 2414 24454 2466 24506
rect 2478 24454 2530 24506
rect 2542 24454 2594 24506
rect 2606 24454 2658 24506
rect 7350 24454 7402 24506
rect 7414 24454 7466 24506
rect 7478 24454 7530 24506
rect 7542 24454 7594 24506
rect 7606 24454 7658 24506
rect 7196 24352 7248 24404
rect 6000 24148 6052 24200
rect 6736 24148 6788 24200
rect 7932 24080 7984 24132
rect 7748 24055 7800 24064
rect 7748 24021 7757 24055
rect 7757 24021 7791 24055
rect 7791 24021 7800 24055
rect 7748 24012 7800 24021
rect 7840 24012 7892 24064
rect 3010 23910 3062 23962
rect 3074 23910 3126 23962
rect 3138 23910 3190 23962
rect 3202 23910 3254 23962
rect 3266 23910 3318 23962
rect 8010 23910 8062 23962
rect 8074 23910 8126 23962
rect 8138 23910 8190 23962
rect 8202 23910 8254 23962
rect 8266 23910 8318 23962
rect 7748 23808 7800 23860
rect 7840 23851 7892 23860
rect 7840 23817 7849 23851
rect 7849 23817 7883 23851
rect 7883 23817 7892 23851
rect 7840 23808 7892 23817
rect 8392 23808 8444 23860
rect 8300 23604 8352 23656
rect 6460 23536 6512 23588
rect 7104 23536 7156 23588
rect 6736 23468 6788 23520
rect 7840 23468 7892 23520
rect 2350 23366 2402 23418
rect 2414 23366 2466 23418
rect 2478 23366 2530 23418
rect 2542 23366 2594 23418
rect 2606 23366 2658 23418
rect 7350 23366 7402 23418
rect 7414 23366 7466 23418
rect 7478 23366 7530 23418
rect 7542 23366 7594 23418
rect 7606 23366 7658 23418
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 6552 23103 6604 23112
rect 6552 23069 6561 23103
rect 6561 23069 6595 23103
rect 6595 23069 6604 23103
rect 6552 23060 6604 23069
rect 6736 22992 6788 23044
rect 6920 22992 6972 23044
rect 7104 22992 7156 23044
rect 3010 22822 3062 22874
rect 3074 22822 3126 22874
rect 3138 22822 3190 22874
rect 3202 22822 3254 22874
rect 3266 22822 3318 22874
rect 8010 22822 8062 22874
rect 8074 22822 8126 22874
rect 8138 22822 8190 22874
rect 8202 22822 8254 22874
rect 8266 22822 8318 22874
rect 7840 22720 7892 22772
rect 8392 22720 8444 22772
rect 7380 22652 7432 22704
rect 7288 22584 7340 22636
rect 7840 22448 7892 22500
rect 7932 22448 7984 22500
rect 6644 22380 6696 22432
rect 7012 22380 7064 22432
rect 7288 22380 7340 22432
rect 7748 22380 7800 22432
rect 2350 22278 2402 22330
rect 2414 22278 2466 22330
rect 2478 22278 2530 22330
rect 2542 22278 2594 22330
rect 2606 22278 2658 22330
rect 7350 22278 7402 22330
rect 7414 22278 7466 22330
rect 7478 22278 7530 22330
rect 7542 22278 7594 22330
rect 7606 22278 7658 22330
rect 6552 22040 6604 22092
rect 6920 21972 6972 22024
rect 7748 21904 7800 21956
rect 7012 21836 7064 21888
rect 3010 21734 3062 21786
rect 3074 21734 3126 21786
rect 3138 21734 3190 21786
rect 3202 21734 3254 21786
rect 3266 21734 3318 21786
rect 8010 21734 8062 21786
rect 8074 21734 8126 21786
rect 8138 21734 8190 21786
rect 8202 21734 8254 21786
rect 8266 21734 8318 21786
rect 8300 21564 8352 21616
rect 7012 21539 7064 21548
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 7932 21428 7984 21480
rect 7748 21335 7800 21344
rect 7748 21301 7757 21335
rect 7757 21301 7791 21335
rect 7791 21301 7800 21335
rect 7748 21292 7800 21301
rect 2350 21190 2402 21242
rect 2414 21190 2466 21242
rect 2478 21190 2530 21242
rect 2542 21190 2594 21242
rect 2606 21190 2658 21242
rect 7350 21190 7402 21242
rect 7414 21190 7466 21242
rect 7478 21190 7530 21242
rect 7542 21190 7594 21242
rect 7606 21190 7658 21242
rect 6920 21088 6972 21140
rect 7288 21088 7340 21140
rect 6552 20995 6604 21004
rect 6552 20961 6561 20995
rect 6561 20961 6595 20995
rect 6595 20961 6604 20995
rect 6552 20952 6604 20961
rect 7104 20816 7156 20868
rect 7288 20816 7340 20868
rect 8392 20748 8444 20800
rect 3010 20646 3062 20698
rect 3074 20646 3126 20698
rect 3138 20646 3190 20698
rect 3202 20646 3254 20698
rect 3266 20646 3318 20698
rect 8010 20646 8062 20698
rect 8074 20646 8126 20698
rect 8138 20646 8190 20698
rect 8202 20646 8254 20698
rect 8266 20646 8318 20698
rect 7104 20544 7156 20596
rect 7748 20544 7800 20596
rect 7932 20544 7984 20596
rect 8208 20476 8260 20528
rect 7932 20408 7984 20460
rect 8116 20451 8168 20460
rect 8116 20417 8125 20451
rect 8125 20417 8159 20451
rect 8159 20417 8168 20451
rect 8116 20408 8168 20417
rect 7196 20340 7248 20392
rect 7840 20272 7892 20324
rect 7104 20204 7156 20256
rect 7288 20204 7340 20256
rect 7748 20247 7800 20256
rect 7748 20213 7757 20247
rect 7757 20213 7791 20247
rect 7791 20213 7800 20247
rect 7748 20204 7800 20213
rect 2350 20102 2402 20154
rect 2414 20102 2466 20154
rect 2478 20102 2530 20154
rect 2542 20102 2594 20154
rect 2606 20102 2658 20154
rect 7350 20102 7402 20154
rect 7414 20102 7466 20154
rect 7478 20102 7530 20154
rect 7542 20102 7594 20154
rect 7606 20102 7658 20154
rect 7748 20000 7800 20052
rect 8116 20000 8168 20052
rect 6736 19932 6788 19984
rect 8392 19907 8444 19916
rect 8392 19873 8401 19907
rect 8401 19873 8435 19907
rect 8435 19873 8444 19907
rect 8392 19864 8444 19873
rect 8300 19728 8352 19780
rect 7196 19660 7248 19712
rect 7840 19660 7892 19712
rect 8208 19660 8260 19712
rect 8392 19660 8444 19712
rect 3010 19558 3062 19610
rect 3074 19558 3126 19610
rect 3138 19558 3190 19610
rect 3202 19558 3254 19610
rect 3266 19558 3318 19610
rect 8010 19558 8062 19610
rect 8074 19558 8126 19610
rect 8138 19558 8190 19610
rect 8202 19558 8254 19610
rect 8266 19558 8318 19610
rect 7196 19456 7248 19508
rect 6736 19388 6788 19440
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 2350 19014 2402 19066
rect 2414 19014 2466 19066
rect 2478 19014 2530 19066
rect 2542 19014 2594 19066
rect 2606 19014 2658 19066
rect 7350 19014 7402 19066
rect 7414 19014 7466 19066
rect 7478 19014 7530 19066
rect 7542 19014 7594 19066
rect 7606 19014 7658 19066
rect 8208 18912 8260 18964
rect 7932 18844 7984 18896
rect 7748 18776 7800 18828
rect 7196 18615 7248 18624
rect 7196 18581 7205 18615
rect 7205 18581 7239 18615
rect 7239 18581 7248 18615
rect 7196 18572 7248 18581
rect 7840 18708 7892 18760
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 3202 18470 3254 18522
rect 3266 18470 3318 18522
rect 8010 18470 8062 18522
rect 8074 18470 8126 18522
rect 8138 18470 8190 18522
rect 8202 18470 8254 18522
rect 8266 18470 8318 18522
rect 7196 18368 7248 18420
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 7932 18232 7984 18284
rect 7288 18164 7340 18216
rect 8392 18028 8444 18080
rect 2350 17926 2402 17978
rect 2414 17926 2466 17978
rect 2478 17926 2530 17978
rect 2542 17926 2594 17978
rect 2606 17926 2658 17978
rect 7350 17926 7402 17978
rect 7414 17926 7466 17978
rect 7478 17926 7530 17978
rect 7542 17926 7594 17978
rect 7606 17926 7658 17978
rect 7840 17824 7892 17876
rect 6920 17552 6972 17604
rect 8484 17552 8536 17604
rect 7104 17484 7156 17536
rect 7748 17527 7800 17536
rect 7748 17493 7757 17527
rect 7757 17493 7791 17527
rect 7791 17493 7800 17527
rect 7748 17484 7800 17493
rect 7840 17484 7892 17536
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 3202 17382 3254 17434
rect 3266 17382 3318 17434
rect 8010 17382 8062 17434
rect 8074 17382 8126 17434
rect 8138 17382 8190 17434
rect 8202 17382 8254 17434
rect 8266 17382 8318 17434
rect 7748 17280 7800 17332
rect 7840 17323 7892 17332
rect 7840 17289 7849 17323
rect 7849 17289 7883 17323
rect 7883 17289 7892 17323
rect 7840 17280 7892 17289
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 6736 17076 6788 17128
rect 8300 17076 8352 17128
rect 6644 17008 6696 17060
rect 6920 16940 6972 16992
rect 7932 16940 7984 16992
rect 2350 16838 2402 16890
rect 2414 16838 2466 16890
rect 2478 16838 2530 16890
rect 2542 16838 2594 16890
rect 2606 16838 2658 16890
rect 7350 16838 7402 16890
rect 7414 16838 7466 16890
rect 7478 16838 7530 16890
rect 7542 16838 7594 16890
rect 7606 16838 7658 16890
rect 6644 16736 6696 16788
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7840 16464 7892 16516
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 3202 16294 3254 16346
rect 3266 16294 3318 16346
rect 8010 16294 8062 16346
rect 8074 16294 8126 16346
rect 8138 16294 8190 16346
rect 8202 16294 8254 16346
rect 8266 16294 8318 16346
rect 6920 16056 6972 16108
rect 7932 16192 7984 16244
rect 7840 15920 7892 15972
rect 7932 15852 7984 15904
rect 2350 15750 2402 15802
rect 2414 15750 2466 15802
rect 2478 15750 2530 15802
rect 2542 15750 2594 15802
rect 2606 15750 2658 15802
rect 7350 15750 7402 15802
rect 7414 15750 7466 15802
rect 7478 15750 7530 15802
rect 7542 15750 7594 15802
rect 7606 15750 7658 15802
rect 7932 15512 7984 15564
rect 6920 15444 6972 15496
rect 8392 15444 8444 15496
rect 6644 15308 6696 15360
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 3202 15206 3254 15258
rect 3266 15206 3318 15258
rect 8010 15206 8062 15258
rect 8074 15206 8126 15258
rect 8138 15206 8190 15258
rect 8202 15206 8254 15258
rect 8266 15206 8318 15258
rect 6552 15104 6604 15156
rect 6828 15036 6880 15088
rect 8392 15104 8444 15156
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 8852 14832 8904 14884
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 8208 14764 8260 14816
rect 2350 14662 2402 14714
rect 2414 14662 2466 14714
rect 2478 14662 2530 14714
rect 2542 14662 2594 14714
rect 2606 14662 2658 14714
rect 7350 14662 7402 14714
rect 7414 14662 7466 14714
rect 7478 14662 7530 14714
rect 7542 14662 7594 14714
rect 7606 14662 7658 14714
rect 6920 14560 6972 14612
rect 7196 14560 7248 14612
rect 7288 14535 7340 14544
rect 7288 14501 7297 14535
rect 7297 14501 7331 14535
rect 7331 14501 7340 14535
rect 7288 14492 7340 14501
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 6092 14331 6144 14340
rect 6092 14297 6101 14331
rect 6101 14297 6135 14331
rect 6135 14297 6144 14331
rect 6092 14288 6144 14297
rect 6460 14288 6512 14340
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 7840 14220 7892 14272
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 3202 14118 3254 14170
rect 3266 14118 3318 14170
rect 8010 14118 8062 14170
rect 8074 14118 8126 14170
rect 8138 14118 8190 14170
rect 8202 14118 8254 14170
rect 8266 14118 8318 14170
rect 6920 13948 6972 14000
rect 7288 13948 7340 14000
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 7840 13812 7892 13864
rect 2350 13574 2402 13626
rect 2414 13574 2466 13626
rect 2478 13574 2530 13626
rect 2542 13574 2594 13626
rect 2606 13574 2658 13626
rect 7350 13574 7402 13626
rect 7414 13574 7466 13626
rect 7478 13574 7530 13626
rect 7542 13574 7594 13626
rect 7606 13574 7658 13626
rect 7840 13336 7892 13388
rect 8300 13200 8352 13252
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 7840 13132 7892 13184
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 3202 13030 3254 13082
rect 3266 13030 3318 13082
rect 8010 13030 8062 13082
rect 8074 13030 8126 13082
rect 8138 13030 8190 13082
rect 8202 13030 8254 13082
rect 8266 13030 8318 13082
rect 6736 12928 6788 12980
rect 7012 12928 7064 12980
rect 7196 12928 7248 12980
rect 6092 12792 6144 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 8300 12631 8352 12640
rect 8300 12597 8309 12631
rect 8309 12597 8343 12631
rect 8343 12597 8352 12631
rect 8300 12588 8352 12597
rect 2350 12486 2402 12538
rect 2414 12486 2466 12538
rect 2478 12486 2530 12538
rect 2542 12486 2594 12538
rect 2606 12486 2658 12538
rect 7350 12486 7402 12538
rect 7414 12486 7466 12538
rect 7478 12486 7530 12538
rect 7542 12486 7594 12538
rect 7606 12486 7658 12538
rect 7840 12248 7892 12300
rect 8576 12248 8628 12300
rect 7932 12180 7984 12232
rect 6736 12112 6788 12164
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 7840 12044 7892 12096
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 3202 11942 3254 11994
rect 3266 11942 3318 11994
rect 8010 11942 8062 11994
rect 8074 11942 8126 11994
rect 8138 11942 8190 11994
rect 8202 11942 8254 11994
rect 8266 11942 8318 11994
rect 6736 11883 6788 11892
rect 6736 11849 6745 11883
rect 6745 11849 6779 11883
rect 6779 11849 6788 11883
rect 6736 11840 6788 11849
rect 7748 11840 7800 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 8484 11636 8536 11688
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7932 11500 7984 11552
rect 2350 11398 2402 11450
rect 2414 11398 2466 11450
rect 2478 11398 2530 11450
rect 2542 11398 2594 11450
rect 2606 11398 2658 11450
rect 7350 11398 7402 11450
rect 7414 11398 7466 11450
rect 7478 11398 7530 11450
rect 7542 11398 7594 11450
rect 7606 11398 7658 11450
rect 7196 11296 7248 11348
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 6828 11203 6880 11212
rect 6828 11169 6837 11203
rect 6837 11169 6871 11203
rect 6871 11169 6880 11203
rect 6828 11160 6880 11169
rect 7012 10956 7064 11008
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 3202 10854 3254 10906
rect 3266 10854 3318 10906
rect 8010 10854 8062 10906
rect 8074 10854 8126 10906
rect 8138 10854 8190 10906
rect 8202 10854 8254 10906
rect 8266 10854 8318 10906
rect 7932 10752 7984 10804
rect 7748 10548 7800 10600
rect 8576 10548 8628 10600
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 2350 10310 2402 10362
rect 2414 10310 2466 10362
rect 2478 10310 2530 10362
rect 2542 10310 2594 10362
rect 2606 10310 2658 10362
rect 7350 10310 7402 10362
rect 7414 10310 7466 10362
rect 7478 10310 7530 10362
rect 7542 10310 7594 10362
rect 7606 10310 7658 10362
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 7196 10072 7248 10124
rect 7288 9936 7340 9988
rect 7012 9868 7064 9920
rect 8392 9868 8444 9920
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 3202 9766 3254 9818
rect 3266 9766 3318 9818
rect 8010 9766 8062 9818
rect 8074 9766 8126 9818
rect 8138 9766 8190 9818
rect 8202 9766 8254 9818
rect 8266 9766 8318 9818
rect 7012 9528 7064 9580
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 6736 9460 6788 9512
rect 7840 9392 7892 9444
rect 7932 9392 7984 9444
rect 8576 9460 8628 9512
rect 7748 9367 7800 9376
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 2350 9222 2402 9274
rect 2414 9222 2466 9274
rect 2478 9222 2530 9274
rect 2542 9222 2594 9274
rect 2606 9222 2658 9274
rect 7350 9222 7402 9274
rect 7414 9222 7466 9274
rect 7478 9222 7530 9274
rect 7542 9222 7594 9274
rect 7606 9222 7658 9274
rect 6736 9163 6788 9172
rect 6736 9129 6745 9163
rect 6745 9129 6779 9163
rect 6779 9129 6788 9163
rect 6736 9120 6788 9129
rect 7748 9120 7800 9172
rect 8116 9120 8168 9172
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 8300 8916 8352 8968
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 8010 8678 8062 8730
rect 8074 8678 8126 8730
rect 8138 8678 8190 8730
rect 8202 8678 8254 8730
rect 8266 8678 8318 8730
rect 7196 8576 7248 8628
rect 7288 8508 7340 8560
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 5080 8236 5132 8288
rect 2350 8134 2402 8186
rect 2414 8134 2466 8186
rect 2478 8134 2530 8186
rect 2542 8134 2594 8186
rect 2606 8134 2658 8186
rect 7350 8134 7402 8186
rect 7414 8134 7466 8186
rect 7478 8134 7530 8186
rect 7542 8134 7594 8186
rect 7606 8134 7658 8186
rect 4804 7964 4856 8016
rect 6552 7964 6604 8016
rect 3976 7896 4028 7948
rect 4160 7760 4212 7812
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 7932 8032 7984 8084
rect 7840 7896 7892 7948
rect 7196 7828 7248 7880
rect 7380 7828 7432 7880
rect 7748 7828 7800 7880
rect 5356 7760 5408 7812
rect 5724 7760 5776 7812
rect 6920 7760 6972 7812
rect 5540 7692 5592 7744
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 7932 7692 7984 7744
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 8010 7590 8062 7642
rect 8074 7590 8126 7642
rect 8138 7590 8190 7642
rect 8202 7590 8254 7642
rect 8266 7590 8318 7642
rect 4160 7488 4212 7540
rect 4436 7488 4488 7540
rect 5724 7488 5776 7540
rect 4804 7420 4856 7472
rect 7748 7488 7800 7540
rect 7380 7420 7432 7472
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 6000 7284 6052 7336
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 6552 7352 6604 7404
rect 6920 7148 6972 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 2350 7046 2402 7098
rect 2414 7046 2466 7098
rect 2478 7046 2530 7098
rect 2542 7046 2594 7098
rect 2606 7046 2658 7098
rect 7350 7046 7402 7098
rect 7414 7046 7466 7098
rect 7478 7046 7530 7098
rect 7542 7046 7594 7098
rect 7606 7046 7658 7098
rect 3884 6944 3936 6996
rect 5540 6944 5592 6996
rect 6920 6944 6972 6996
rect 7012 6876 7064 6928
rect 7104 6740 7156 6792
rect 3976 6672 4028 6724
rect 4804 6672 4856 6724
rect 5632 6672 5684 6724
rect 7840 6808 7892 6860
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 7840 6604 7892 6656
rect 8484 6604 8536 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 8010 6502 8062 6554
rect 8074 6502 8126 6554
rect 8138 6502 8190 6554
rect 8202 6502 8254 6554
rect 8266 6502 8318 6554
rect 7104 6400 7156 6452
rect 7840 6443 7892 6452
rect 7840 6409 7849 6443
rect 7849 6409 7883 6443
rect 7883 6409 7892 6443
rect 7840 6400 7892 6409
rect 7656 6375 7708 6384
rect 7656 6341 7665 6375
rect 7665 6341 7699 6375
rect 7699 6341 7708 6375
rect 7656 6332 7708 6341
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 2350 5958 2402 6010
rect 2414 5958 2466 6010
rect 2478 5958 2530 6010
rect 2542 5958 2594 6010
rect 2606 5958 2658 6010
rect 7350 5958 7402 6010
rect 7414 5958 7466 6010
rect 7478 5958 7530 6010
rect 7542 5958 7594 6010
rect 7606 5958 7658 6010
rect 8484 5856 8536 5908
rect 8852 5652 8904 5704
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 8010 5414 8062 5466
rect 8074 5414 8126 5466
rect 8138 5414 8190 5466
rect 8202 5414 8254 5466
rect 8266 5414 8318 5466
rect 2350 4870 2402 4922
rect 2414 4870 2466 4922
rect 2478 4870 2530 4922
rect 2542 4870 2594 4922
rect 2606 4870 2658 4922
rect 7350 4870 7402 4922
rect 7414 4870 7466 4922
rect 7478 4870 7530 4922
rect 7542 4870 7594 4922
rect 7606 4870 7658 4922
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 8010 4326 8062 4378
rect 8074 4326 8126 4378
rect 8138 4326 8190 4378
rect 8202 4326 8254 4378
rect 8266 4326 8318 4378
rect 2350 3782 2402 3834
rect 2414 3782 2466 3834
rect 2478 3782 2530 3834
rect 2542 3782 2594 3834
rect 2606 3782 2658 3834
rect 7350 3782 7402 3834
rect 7414 3782 7466 3834
rect 7478 3782 7530 3834
rect 7542 3782 7594 3834
rect 7606 3782 7658 3834
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 8010 3238 8062 3290
rect 8074 3238 8126 3290
rect 8138 3238 8190 3290
rect 8202 3238 8254 3290
rect 8266 3238 8318 3290
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 848 2796 900 2848
rect 2136 2839 2188 2848
rect 2136 2805 2145 2839
rect 2145 2805 2179 2839
rect 2179 2805 2188 2839
rect 2136 2796 2188 2805
rect 2350 2694 2402 2746
rect 2414 2694 2466 2746
rect 2478 2694 2530 2746
rect 2542 2694 2594 2746
rect 2606 2694 2658 2746
rect 7350 2694 7402 2746
rect 7414 2694 7466 2746
rect 7478 2694 7530 2746
rect 7542 2694 7594 2746
rect 7606 2694 7658 2746
rect 7748 2592 7800 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 5540 2388 5592 2440
rect 5816 2388 5868 2440
rect 7656 2363 7708 2372
rect 7656 2329 7665 2363
rect 7665 2329 7699 2363
rect 7699 2329 7708 2363
rect 7656 2320 7708 2329
rect 9128 2320 9180 2372
rect 4160 2295 4212 2304
rect 4160 2261 4169 2295
rect 4169 2261 4203 2295
rect 4203 2261 4212 2295
rect 4160 2252 4212 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 8010 2150 8062 2202
rect 8074 2150 8126 2202
rect 8138 2150 8190 2202
rect 8202 2150 8254 2202
rect 8266 2150 8318 2202
<< metal2 >>
rect 2502 79200 2558 80000
rect 7208 79206 7420 79234
rect 2516 78282 2544 79200
rect 2516 78254 2728 78282
rect 2350 77820 2658 77829
rect 2350 77818 2356 77820
rect 2412 77818 2436 77820
rect 2492 77818 2516 77820
rect 2572 77818 2596 77820
rect 2652 77818 2658 77820
rect 2412 77766 2414 77818
rect 2594 77766 2596 77818
rect 2350 77764 2356 77766
rect 2412 77764 2436 77766
rect 2492 77764 2516 77766
rect 2572 77764 2596 77766
rect 2652 77764 2658 77766
rect 2350 77755 2658 77764
rect 2700 77518 2728 78254
rect 2688 77512 2740 77518
rect 2688 77454 2740 77460
rect 5540 77444 5592 77450
rect 5540 77386 5592 77392
rect 3010 77276 3318 77285
rect 3010 77274 3016 77276
rect 3072 77274 3096 77276
rect 3152 77274 3176 77276
rect 3232 77274 3256 77276
rect 3312 77274 3318 77276
rect 3072 77222 3074 77274
rect 3254 77222 3256 77274
rect 3010 77220 3016 77222
rect 3072 77220 3096 77222
rect 3152 77220 3176 77222
rect 3232 77220 3256 77222
rect 3312 77220 3318 77222
rect 3010 77211 3318 77220
rect 2350 76732 2658 76741
rect 2350 76730 2356 76732
rect 2412 76730 2436 76732
rect 2492 76730 2516 76732
rect 2572 76730 2596 76732
rect 2652 76730 2658 76732
rect 2412 76678 2414 76730
rect 2594 76678 2596 76730
rect 2350 76676 2356 76678
rect 2412 76676 2436 76678
rect 2492 76676 2516 76678
rect 2572 76676 2596 76678
rect 2652 76676 2658 76678
rect 2350 76667 2658 76676
rect 3010 76188 3318 76197
rect 3010 76186 3016 76188
rect 3072 76186 3096 76188
rect 3152 76186 3176 76188
rect 3232 76186 3256 76188
rect 3312 76186 3318 76188
rect 3072 76134 3074 76186
rect 3254 76134 3256 76186
rect 3010 76132 3016 76134
rect 3072 76132 3096 76134
rect 3152 76132 3176 76134
rect 3232 76132 3256 76134
rect 3312 76132 3318 76134
rect 3010 76123 3318 76132
rect 2350 75644 2658 75653
rect 2350 75642 2356 75644
rect 2412 75642 2436 75644
rect 2492 75642 2516 75644
rect 2572 75642 2596 75644
rect 2652 75642 2658 75644
rect 2412 75590 2414 75642
rect 2594 75590 2596 75642
rect 2350 75588 2356 75590
rect 2412 75588 2436 75590
rect 2492 75588 2516 75590
rect 2572 75588 2596 75590
rect 2652 75588 2658 75590
rect 2350 75579 2658 75588
rect 3010 75100 3318 75109
rect 3010 75098 3016 75100
rect 3072 75098 3096 75100
rect 3152 75098 3176 75100
rect 3232 75098 3256 75100
rect 3312 75098 3318 75100
rect 3072 75046 3074 75098
rect 3254 75046 3256 75098
rect 3010 75044 3016 75046
rect 3072 75044 3096 75046
rect 3152 75044 3176 75046
rect 3232 75044 3256 75046
rect 3312 75044 3318 75046
rect 3010 75035 3318 75044
rect 2350 74556 2658 74565
rect 2350 74554 2356 74556
rect 2412 74554 2436 74556
rect 2492 74554 2516 74556
rect 2572 74554 2596 74556
rect 2652 74554 2658 74556
rect 2412 74502 2414 74554
rect 2594 74502 2596 74554
rect 2350 74500 2356 74502
rect 2412 74500 2436 74502
rect 2492 74500 2516 74502
rect 2572 74500 2596 74502
rect 2652 74500 2658 74502
rect 2350 74491 2658 74500
rect 3010 74012 3318 74021
rect 3010 74010 3016 74012
rect 3072 74010 3096 74012
rect 3152 74010 3176 74012
rect 3232 74010 3256 74012
rect 3312 74010 3318 74012
rect 3072 73958 3074 74010
rect 3254 73958 3256 74010
rect 3010 73956 3016 73958
rect 3072 73956 3096 73958
rect 3152 73956 3176 73958
rect 3232 73956 3256 73958
rect 3312 73956 3318 73958
rect 3010 73947 3318 73956
rect 5552 73778 5580 77386
rect 5540 73772 5592 73778
rect 5540 73714 5592 73720
rect 6368 73772 6420 73778
rect 6368 73714 6420 73720
rect 2350 73468 2658 73477
rect 2350 73466 2356 73468
rect 2412 73466 2436 73468
rect 2492 73466 2516 73468
rect 2572 73466 2596 73468
rect 2652 73466 2658 73468
rect 2412 73414 2414 73466
rect 2594 73414 2596 73466
rect 2350 73412 2356 73414
rect 2412 73412 2436 73414
rect 2492 73412 2516 73414
rect 2572 73412 2596 73414
rect 2652 73412 2658 73414
rect 2350 73403 2658 73412
rect 5080 73160 5132 73166
rect 5080 73102 5132 73108
rect 3010 72924 3318 72933
rect 3010 72922 3016 72924
rect 3072 72922 3096 72924
rect 3152 72922 3176 72924
rect 3232 72922 3256 72924
rect 3312 72922 3318 72924
rect 3072 72870 3074 72922
rect 3254 72870 3256 72922
rect 3010 72868 3016 72870
rect 3072 72868 3096 72870
rect 3152 72868 3176 72870
rect 3232 72868 3256 72870
rect 3312 72868 3318 72870
rect 3010 72859 3318 72868
rect 2350 72380 2658 72389
rect 2350 72378 2356 72380
rect 2412 72378 2436 72380
rect 2492 72378 2516 72380
rect 2572 72378 2596 72380
rect 2652 72378 2658 72380
rect 2412 72326 2414 72378
rect 2594 72326 2596 72378
rect 2350 72324 2356 72326
rect 2412 72324 2436 72326
rect 2492 72324 2516 72326
rect 2572 72324 2596 72326
rect 2652 72324 2658 72326
rect 2350 72315 2658 72324
rect 5092 72146 5120 73102
rect 5356 73092 5408 73098
rect 5356 73034 5408 73040
rect 5368 72826 5396 73034
rect 5356 72820 5408 72826
rect 5356 72762 5408 72768
rect 4436 72140 4488 72146
rect 4436 72082 4488 72088
rect 5080 72140 5132 72146
rect 5080 72082 5132 72088
rect 3010 71836 3318 71845
rect 3010 71834 3016 71836
rect 3072 71834 3096 71836
rect 3152 71834 3176 71836
rect 3232 71834 3256 71836
rect 3312 71834 3318 71836
rect 3072 71782 3074 71834
rect 3254 71782 3256 71834
rect 3010 71780 3016 71782
rect 3072 71780 3096 71782
rect 3152 71780 3176 71782
rect 3232 71780 3256 71782
rect 3312 71780 3318 71782
rect 3010 71771 3318 71780
rect 2350 71292 2658 71301
rect 2350 71290 2356 71292
rect 2412 71290 2436 71292
rect 2492 71290 2516 71292
rect 2572 71290 2596 71292
rect 2652 71290 2658 71292
rect 2412 71238 2414 71290
rect 2594 71238 2596 71290
rect 2350 71236 2356 71238
rect 2412 71236 2436 71238
rect 2492 71236 2516 71238
rect 2572 71236 2596 71238
rect 2652 71236 2658 71238
rect 2350 71227 2658 71236
rect 3010 70748 3318 70757
rect 3010 70746 3016 70748
rect 3072 70746 3096 70748
rect 3152 70746 3176 70748
rect 3232 70746 3256 70748
rect 3312 70746 3318 70748
rect 3072 70694 3074 70746
rect 3254 70694 3256 70746
rect 3010 70692 3016 70694
rect 3072 70692 3096 70694
rect 3152 70692 3176 70694
rect 3232 70692 3256 70694
rect 3312 70692 3318 70694
rect 3010 70683 3318 70692
rect 4448 70514 4476 72082
rect 5080 72004 5132 72010
rect 5080 71946 5132 71952
rect 5092 71738 5120 71946
rect 5816 71936 5868 71942
rect 5816 71878 5868 71884
rect 5080 71732 5132 71738
rect 5080 71674 5132 71680
rect 4988 70848 5040 70854
rect 4988 70790 5040 70796
rect 5000 70582 5028 70790
rect 4988 70576 5040 70582
rect 4988 70518 5040 70524
rect 5828 70514 5856 71878
rect 5908 71528 5960 71534
rect 5908 71470 5960 71476
rect 5920 70990 5948 71470
rect 6092 71392 6144 71398
rect 6092 71334 6144 71340
rect 6104 71058 6132 71334
rect 6092 71052 6144 71058
rect 6092 70994 6144 71000
rect 5908 70984 5960 70990
rect 5908 70926 5960 70932
rect 4436 70508 4488 70514
rect 4436 70450 4488 70456
rect 5816 70508 5868 70514
rect 5816 70450 5868 70456
rect 2350 70204 2658 70213
rect 2350 70202 2356 70204
rect 2412 70202 2436 70204
rect 2492 70202 2516 70204
rect 2572 70202 2596 70204
rect 2652 70202 2658 70204
rect 2412 70150 2414 70202
rect 2594 70150 2596 70202
rect 2350 70148 2356 70150
rect 2412 70148 2436 70150
rect 2492 70148 2516 70150
rect 2572 70148 2596 70150
rect 2652 70148 2658 70150
rect 2350 70139 2658 70148
rect 3010 69660 3318 69669
rect 3010 69658 3016 69660
rect 3072 69658 3096 69660
rect 3152 69658 3176 69660
rect 3232 69658 3256 69660
rect 3312 69658 3318 69660
rect 3072 69606 3074 69658
rect 3254 69606 3256 69658
rect 3010 69604 3016 69606
rect 3072 69604 3096 69606
rect 3152 69604 3176 69606
rect 3232 69604 3256 69606
rect 3312 69604 3318 69606
rect 3010 69595 3318 69604
rect 4448 69426 4476 70450
rect 5908 69760 5960 69766
rect 5908 69702 5960 69708
rect 4436 69420 4488 69426
rect 4436 69362 4488 69368
rect 2350 69116 2658 69125
rect 2350 69114 2356 69116
rect 2412 69114 2436 69116
rect 2492 69114 2516 69116
rect 2572 69114 2596 69116
rect 2652 69114 2658 69116
rect 2412 69062 2414 69114
rect 2594 69062 2596 69114
rect 2350 69060 2356 69062
rect 2412 69060 2436 69062
rect 2492 69060 2516 69062
rect 2572 69060 2596 69062
rect 2652 69060 2658 69062
rect 2350 69051 2658 69060
rect 3010 68572 3318 68581
rect 3010 68570 3016 68572
rect 3072 68570 3096 68572
rect 3152 68570 3176 68572
rect 3232 68570 3256 68572
rect 3312 68570 3318 68572
rect 3072 68518 3074 68570
rect 3254 68518 3256 68570
rect 3010 68516 3016 68518
rect 3072 68516 3096 68518
rect 3152 68516 3176 68518
rect 3232 68516 3256 68518
rect 3312 68516 3318 68518
rect 3010 68507 3318 68516
rect 2350 68028 2658 68037
rect 2350 68026 2356 68028
rect 2412 68026 2436 68028
rect 2492 68026 2516 68028
rect 2572 68026 2596 68028
rect 2652 68026 2658 68028
rect 2412 67974 2414 68026
rect 2594 67974 2596 68026
rect 2350 67972 2356 67974
rect 2412 67972 2436 67974
rect 2492 67972 2516 67974
rect 2572 67972 2596 67974
rect 2652 67972 2658 67974
rect 2350 67963 2658 67972
rect 4448 67794 4476 69362
rect 4712 69352 4764 69358
rect 4712 69294 4764 69300
rect 4724 69018 4752 69294
rect 4712 69012 4764 69018
rect 4712 68954 4764 68960
rect 5920 68814 5948 69702
rect 6104 69578 6132 70994
rect 6184 70848 6236 70854
rect 6184 70790 6236 70796
rect 6196 70446 6224 70790
rect 6184 70440 6236 70446
rect 6184 70382 6236 70388
rect 6380 70394 6408 73714
rect 6736 73704 6788 73710
rect 6736 73646 6788 73652
rect 7012 73704 7064 73710
rect 7012 73646 7064 73652
rect 6644 73568 6696 73574
rect 6644 73510 6696 73516
rect 6656 73098 6684 73510
rect 6644 73092 6696 73098
rect 6644 73034 6696 73040
rect 6656 72842 6684 73034
rect 6564 72826 6684 72842
rect 6564 72820 6696 72826
rect 6564 72814 6644 72820
rect 6460 72480 6512 72486
rect 6460 72422 6512 72428
rect 6472 71466 6500 72422
rect 6564 72078 6592 72814
rect 6644 72762 6696 72768
rect 6644 72684 6696 72690
rect 6644 72626 6696 72632
rect 6552 72072 6604 72078
rect 6552 72014 6604 72020
rect 6552 71936 6604 71942
rect 6552 71878 6604 71884
rect 6564 71534 6592 71878
rect 6552 71528 6604 71534
rect 6552 71470 6604 71476
rect 6460 71460 6512 71466
rect 6460 71402 6512 71408
rect 6656 70394 6684 72626
rect 6748 72146 6776 73646
rect 7024 73370 7052 73646
rect 7012 73364 7064 73370
rect 7012 73306 7064 73312
rect 6828 73024 6880 73030
rect 6828 72966 6880 72972
rect 6840 72622 6868 72966
rect 7012 72684 7064 72690
rect 7012 72626 7064 72632
rect 6828 72616 6880 72622
rect 6828 72558 6880 72564
rect 6736 72140 6788 72146
rect 6736 72082 6788 72088
rect 6748 70514 6776 72082
rect 6840 71738 6868 72558
rect 7024 71738 7052 72626
rect 7104 72480 7156 72486
rect 7104 72422 7156 72428
rect 7116 72146 7144 72422
rect 7104 72140 7156 72146
rect 7104 72082 7156 72088
rect 7104 72004 7156 72010
rect 7104 71946 7156 71952
rect 6828 71732 6880 71738
rect 6828 71674 6880 71680
rect 7012 71732 7064 71738
rect 7012 71674 7064 71680
rect 6920 70984 6972 70990
rect 6920 70926 6972 70932
rect 6736 70508 6788 70514
rect 6736 70450 6788 70456
rect 6196 69766 6224 70382
rect 6380 70366 6500 70394
rect 6184 69760 6236 69766
rect 6184 69702 6236 69708
rect 6104 69550 6316 69578
rect 6000 69352 6052 69358
rect 6000 69294 6052 69300
rect 6012 68882 6040 69294
rect 6288 68882 6316 69550
rect 6000 68876 6052 68882
rect 6000 68818 6052 68824
rect 6276 68876 6328 68882
rect 6276 68818 6328 68824
rect 5908 68808 5960 68814
rect 5908 68750 5960 68756
rect 6012 68474 6040 68818
rect 6000 68468 6052 68474
rect 6000 68410 6052 68416
rect 5172 68128 5224 68134
rect 5172 68070 5224 68076
rect 5184 67794 5212 68070
rect 4436 67788 4488 67794
rect 4436 67730 4488 67736
rect 5172 67788 5224 67794
rect 5172 67730 5224 67736
rect 3010 67484 3318 67493
rect 3010 67482 3016 67484
rect 3072 67482 3096 67484
rect 3152 67482 3176 67484
rect 3232 67482 3256 67484
rect 3312 67482 3318 67484
rect 3072 67430 3074 67482
rect 3254 67430 3256 67482
rect 3010 67428 3016 67430
rect 3072 67428 3096 67430
rect 3152 67428 3176 67430
rect 3232 67428 3256 67430
rect 3312 67428 3318 67430
rect 3010 67419 3318 67428
rect 2350 66940 2658 66949
rect 2350 66938 2356 66940
rect 2412 66938 2436 66940
rect 2492 66938 2516 66940
rect 2572 66938 2596 66940
rect 2652 66938 2658 66940
rect 2412 66886 2414 66938
rect 2594 66886 2596 66938
rect 2350 66884 2356 66886
rect 2412 66884 2436 66886
rect 2492 66884 2516 66886
rect 2572 66884 2596 66886
rect 2652 66884 2658 66886
rect 2350 66875 2658 66884
rect 4448 66706 4476 67730
rect 6092 67584 6144 67590
rect 6092 67526 6144 67532
rect 4436 66700 4488 66706
rect 4436 66642 4488 66648
rect 3010 66396 3318 66405
rect 3010 66394 3016 66396
rect 3072 66394 3096 66396
rect 3152 66394 3176 66396
rect 3232 66394 3256 66396
rect 3312 66394 3318 66396
rect 3072 66342 3074 66394
rect 3254 66342 3256 66394
rect 3010 66340 3016 66342
rect 3072 66340 3096 66342
rect 3152 66340 3176 66342
rect 3232 66340 3256 66342
rect 3312 66340 3318 66342
rect 3010 66331 3318 66340
rect 2350 65852 2658 65861
rect 2350 65850 2356 65852
rect 2412 65850 2436 65852
rect 2492 65850 2516 65852
rect 2572 65850 2596 65852
rect 2652 65850 2658 65852
rect 2412 65798 2414 65850
rect 2594 65798 2596 65850
rect 2350 65796 2356 65798
rect 2412 65796 2436 65798
rect 2492 65796 2516 65798
rect 2572 65796 2596 65798
rect 2652 65796 2658 65798
rect 2350 65787 2658 65796
rect 4448 65618 4476 66642
rect 6104 66638 6132 67526
rect 6092 66632 6144 66638
rect 6092 66574 6144 66580
rect 5080 66564 5132 66570
rect 5080 66506 5132 66512
rect 5092 66298 5120 66506
rect 5724 66496 5776 66502
rect 5724 66438 5776 66444
rect 5080 66292 5132 66298
rect 5080 66234 5132 66240
rect 4436 65612 4488 65618
rect 4436 65554 4488 65560
rect 3010 65308 3318 65317
rect 3010 65306 3016 65308
rect 3072 65306 3096 65308
rect 3152 65306 3176 65308
rect 3232 65306 3256 65308
rect 3312 65306 3318 65308
rect 3072 65254 3074 65306
rect 3254 65254 3256 65306
rect 3010 65252 3016 65254
rect 3072 65252 3096 65254
rect 3152 65252 3176 65254
rect 3232 65252 3256 65254
rect 3312 65252 3318 65254
rect 3010 65243 3318 65252
rect 4448 65142 4476 65554
rect 5080 65476 5132 65482
rect 5080 65418 5132 65424
rect 5092 65210 5120 65418
rect 5736 65362 5764 66438
rect 5816 65612 5868 65618
rect 5816 65554 5868 65560
rect 5552 65334 5764 65362
rect 5080 65204 5132 65210
rect 5080 65146 5132 65152
rect 4436 65136 4488 65142
rect 4356 65084 4436 65090
rect 4356 65078 4488 65084
rect 4356 65062 4476 65078
rect 5552 65074 5580 65334
rect 5540 65068 5592 65074
rect 2350 64764 2658 64773
rect 2350 64762 2356 64764
rect 2412 64762 2436 64764
rect 2492 64762 2516 64764
rect 2572 64762 2596 64764
rect 2652 64762 2658 64764
rect 2412 64710 2414 64762
rect 2594 64710 2596 64762
rect 2350 64708 2356 64710
rect 2412 64708 2436 64710
rect 2492 64708 2516 64710
rect 2572 64708 2596 64710
rect 2652 64708 2658 64710
rect 2350 64699 2658 64708
rect 3010 64220 3318 64229
rect 3010 64218 3016 64220
rect 3072 64218 3096 64220
rect 3152 64218 3176 64220
rect 3232 64218 3256 64220
rect 3312 64218 3318 64220
rect 3072 64166 3074 64218
rect 3254 64166 3256 64218
rect 3010 64164 3016 64166
rect 3072 64164 3096 64166
rect 3152 64164 3176 64166
rect 3232 64164 3256 64166
rect 3312 64164 3318 64166
rect 3010 64155 3318 64164
rect 2350 63676 2658 63685
rect 2350 63674 2356 63676
rect 2412 63674 2436 63676
rect 2492 63674 2516 63676
rect 2572 63674 2596 63676
rect 2652 63674 2658 63676
rect 2412 63622 2414 63674
rect 2594 63622 2596 63674
rect 2350 63620 2356 63622
rect 2412 63620 2436 63622
rect 2492 63620 2516 63622
rect 2572 63620 2596 63622
rect 2652 63620 2658 63622
rect 2350 63611 2658 63620
rect 4356 63442 4384 65062
rect 5540 65010 5592 65016
rect 4804 63776 4856 63782
rect 4804 63718 4856 63724
rect 4816 63578 4844 63718
rect 4804 63572 4856 63578
rect 4804 63514 4856 63520
rect 4344 63436 4396 63442
rect 4344 63378 4396 63384
rect 3010 63132 3318 63141
rect 3010 63130 3016 63132
rect 3072 63130 3096 63132
rect 3152 63130 3176 63132
rect 3232 63130 3256 63132
rect 3312 63130 3318 63132
rect 3072 63078 3074 63130
rect 3254 63078 3256 63130
rect 3010 63076 3016 63078
rect 3072 63076 3096 63078
rect 3152 63076 3176 63078
rect 3232 63076 3256 63078
rect 3312 63076 3318 63078
rect 3010 63067 3318 63076
rect 2350 62588 2658 62597
rect 2350 62586 2356 62588
rect 2412 62586 2436 62588
rect 2492 62586 2516 62588
rect 2572 62586 2596 62588
rect 2652 62586 2658 62588
rect 2412 62534 2414 62586
rect 2594 62534 2596 62586
rect 2350 62532 2356 62534
rect 2412 62532 2436 62534
rect 2492 62532 2516 62534
rect 2572 62532 2596 62534
rect 2652 62532 2658 62534
rect 2350 62523 2658 62532
rect 4356 62354 4384 63378
rect 4712 62688 4764 62694
rect 4712 62630 4764 62636
rect 4724 62354 4752 62630
rect 4344 62348 4396 62354
rect 4344 62290 4396 62296
rect 4712 62348 4764 62354
rect 4712 62290 4764 62296
rect 3010 62044 3318 62053
rect 3010 62042 3016 62044
rect 3072 62042 3096 62044
rect 3152 62042 3176 62044
rect 3232 62042 3256 62044
rect 3312 62042 3318 62044
rect 3072 61990 3074 62042
rect 3254 61990 3256 62042
rect 3010 61988 3016 61990
rect 3072 61988 3096 61990
rect 3152 61988 3176 61990
rect 3232 61988 3256 61990
rect 3312 61988 3318 61990
rect 3010 61979 3318 61988
rect 2350 61500 2658 61509
rect 2350 61498 2356 61500
rect 2412 61498 2436 61500
rect 2492 61498 2516 61500
rect 2572 61498 2596 61500
rect 2652 61498 2658 61500
rect 2412 61446 2414 61498
rect 2594 61446 2596 61498
rect 2350 61444 2356 61446
rect 2412 61444 2436 61446
rect 2492 61444 2516 61446
rect 2572 61444 2596 61446
rect 2652 61444 2658 61446
rect 2350 61435 2658 61444
rect 4356 61266 4384 62290
rect 4344 61260 4396 61266
rect 4344 61202 4396 61208
rect 3010 60956 3318 60965
rect 3010 60954 3016 60956
rect 3072 60954 3096 60956
rect 3152 60954 3176 60956
rect 3232 60954 3256 60956
rect 3312 60954 3318 60956
rect 3072 60902 3074 60954
rect 3254 60902 3256 60954
rect 3010 60900 3016 60902
rect 3072 60900 3096 60902
rect 3152 60900 3176 60902
rect 3232 60900 3256 60902
rect 3312 60900 3318 60902
rect 3010 60891 3318 60900
rect 4356 60734 4384 61202
rect 4712 61124 4764 61130
rect 4712 61066 4764 61072
rect 4724 60858 4752 61066
rect 4712 60852 4764 60858
rect 4712 60794 4764 60800
rect 4356 60706 4476 60734
rect 2350 60412 2658 60421
rect 2350 60410 2356 60412
rect 2412 60410 2436 60412
rect 2492 60410 2516 60412
rect 2572 60410 2596 60412
rect 2652 60410 2658 60412
rect 2412 60358 2414 60410
rect 2594 60358 2596 60410
rect 2350 60356 2356 60358
rect 2412 60356 2436 60358
rect 2492 60356 2516 60358
rect 2572 60356 2596 60358
rect 2652 60356 2658 60358
rect 2350 60347 2658 60356
rect 3010 59868 3318 59877
rect 3010 59866 3016 59868
rect 3072 59866 3096 59868
rect 3152 59866 3176 59868
rect 3232 59866 3256 59868
rect 3312 59866 3318 59868
rect 3072 59814 3074 59866
rect 3254 59814 3256 59866
rect 3010 59812 3016 59814
rect 3072 59812 3096 59814
rect 3152 59812 3176 59814
rect 3232 59812 3256 59814
rect 3312 59812 3318 59814
rect 3010 59803 3318 59812
rect 4448 59634 4476 60706
rect 4896 59968 4948 59974
rect 4896 59910 4948 59916
rect 4908 59770 4936 59910
rect 4896 59764 4948 59770
rect 4896 59706 4948 59712
rect 4436 59628 4488 59634
rect 4436 59570 4488 59576
rect 2350 59324 2658 59333
rect 2350 59322 2356 59324
rect 2412 59322 2436 59324
rect 2492 59322 2516 59324
rect 2572 59322 2596 59324
rect 2652 59322 2658 59324
rect 2412 59270 2414 59322
rect 2594 59270 2596 59322
rect 2350 59268 2356 59270
rect 2412 59268 2436 59270
rect 2492 59268 2516 59270
rect 2572 59268 2596 59270
rect 2652 59268 2658 59270
rect 2350 59259 2658 59268
rect 5264 58880 5316 58886
rect 5264 58822 5316 58828
rect 3010 58780 3318 58789
rect 3010 58778 3016 58780
rect 3072 58778 3096 58780
rect 3152 58778 3176 58780
rect 3232 58778 3256 58780
rect 3312 58778 3318 58780
rect 3072 58726 3074 58778
rect 3254 58726 3256 58778
rect 3010 58724 3016 58726
rect 3072 58724 3096 58726
rect 3152 58724 3176 58726
rect 3232 58724 3256 58726
rect 3312 58724 3318 58726
rect 3010 58715 3318 58724
rect 4712 58608 4764 58614
rect 4712 58550 4764 58556
rect 2350 58236 2658 58245
rect 2350 58234 2356 58236
rect 2412 58234 2436 58236
rect 2492 58234 2516 58236
rect 2572 58234 2596 58236
rect 2652 58234 2658 58236
rect 2412 58182 2414 58234
rect 2594 58182 2596 58234
rect 2350 58180 2356 58182
rect 2412 58180 2436 58182
rect 2492 58180 2516 58182
rect 2572 58180 2596 58182
rect 2652 58180 2658 58182
rect 2350 58171 2658 58180
rect 4724 58138 4752 58550
rect 4712 58132 4764 58138
rect 4712 58074 4764 58080
rect 5276 57934 5304 58822
rect 5264 57928 5316 57934
rect 5264 57870 5316 57876
rect 3010 57692 3318 57701
rect 3010 57690 3016 57692
rect 3072 57690 3096 57692
rect 3152 57690 3176 57692
rect 3232 57690 3256 57692
rect 3312 57690 3318 57692
rect 3072 57638 3074 57690
rect 3254 57638 3256 57690
rect 3010 57636 3016 57638
rect 3072 57636 3096 57638
rect 3152 57636 3176 57638
rect 3232 57636 3256 57638
rect 3312 57636 3318 57638
rect 3010 57627 3318 57636
rect 4712 57384 4764 57390
rect 4712 57326 4764 57332
rect 2350 57148 2658 57157
rect 2350 57146 2356 57148
rect 2412 57146 2436 57148
rect 2492 57146 2516 57148
rect 2572 57146 2596 57148
rect 2652 57146 2658 57148
rect 2412 57094 2414 57146
rect 2594 57094 2596 57146
rect 2350 57092 2356 57094
rect 2412 57092 2436 57094
rect 2492 57092 2516 57094
rect 2572 57092 2596 57094
rect 2652 57092 2658 57094
rect 2350 57083 2658 57092
rect 4724 57050 4752 57326
rect 4712 57044 4764 57050
rect 4712 56986 4764 56992
rect 3010 56604 3318 56613
rect 3010 56602 3016 56604
rect 3072 56602 3096 56604
rect 3152 56602 3176 56604
rect 3232 56602 3256 56604
rect 3312 56602 3318 56604
rect 3072 56550 3074 56602
rect 3254 56550 3256 56602
rect 3010 56548 3016 56550
rect 3072 56548 3096 56550
rect 3152 56548 3176 56550
rect 3232 56548 3256 56550
rect 3312 56548 3318 56550
rect 3010 56539 3318 56548
rect 4896 56160 4948 56166
rect 4896 56102 4948 56108
rect 2350 56060 2658 56069
rect 2350 56058 2356 56060
rect 2412 56058 2436 56060
rect 2492 56058 2516 56060
rect 2572 56058 2596 56060
rect 2652 56058 2658 56060
rect 2412 56006 2414 56058
rect 2594 56006 2596 56058
rect 2350 56004 2356 56006
rect 2412 56004 2436 56006
rect 2492 56004 2516 56006
rect 2572 56004 2596 56006
rect 2652 56004 2658 56006
rect 2350 55995 2658 56004
rect 4908 55826 4936 56102
rect 4896 55820 4948 55826
rect 4896 55762 4948 55768
rect 4436 55752 4488 55758
rect 4436 55694 4488 55700
rect 3010 55516 3318 55525
rect 3010 55514 3016 55516
rect 3072 55514 3096 55516
rect 3152 55514 3176 55516
rect 3232 55514 3256 55516
rect 3312 55514 3318 55516
rect 3072 55462 3074 55514
rect 3254 55462 3256 55514
rect 3010 55460 3016 55462
rect 3072 55460 3096 55462
rect 3152 55460 3176 55462
rect 3232 55460 3256 55462
rect 3312 55460 3318 55462
rect 3010 55451 3318 55460
rect 2350 54972 2658 54981
rect 2350 54970 2356 54972
rect 2412 54970 2436 54972
rect 2492 54970 2516 54972
rect 2572 54970 2596 54972
rect 2652 54970 2658 54972
rect 2412 54918 2414 54970
rect 2594 54918 2596 54970
rect 2350 54916 2356 54918
rect 2412 54916 2436 54918
rect 2492 54916 2516 54918
rect 2572 54916 2596 54918
rect 2652 54916 2658 54918
rect 2350 54907 2658 54916
rect 4448 54670 4476 55694
rect 4436 54664 4488 54670
rect 4436 54606 4488 54612
rect 3010 54428 3318 54437
rect 3010 54426 3016 54428
rect 3072 54426 3096 54428
rect 3152 54426 3176 54428
rect 3232 54426 3256 54428
rect 3312 54426 3318 54428
rect 3072 54374 3074 54426
rect 3254 54374 3256 54426
rect 3010 54372 3016 54374
rect 3072 54372 3096 54374
rect 3152 54372 3176 54374
rect 3232 54372 3256 54374
rect 3312 54372 3318 54374
rect 3010 54363 3318 54372
rect 2350 53884 2658 53893
rect 2350 53882 2356 53884
rect 2412 53882 2436 53884
rect 2492 53882 2516 53884
rect 2572 53882 2596 53884
rect 2652 53882 2658 53884
rect 2412 53830 2414 53882
rect 2594 53830 2596 53882
rect 2350 53828 2356 53830
rect 2412 53828 2436 53830
rect 2492 53828 2516 53830
rect 2572 53828 2596 53830
rect 2652 53828 2658 53830
rect 2350 53819 2658 53828
rect 3010 53340 3318 53349
rect 3010 53338 3016 53340
rect 3072 53338 3096 53340
rect 3152 53338 3176 53340
rect 3232 53338 3256 53340
rect 3312 53338 3318 53340
rect 3072 53286 3074 53338
rect 3254 53286 3256 53338
rect 3010 53284 3016 53286
rect 3072 53284 3096 53286
rect 3152 53284 3176 53286
rect 3232 53284 3256 53286
rect 3312 53284 3318 53286
rect 3010 53275 3318 53284
rect 4448 53038 4476 54606
rect 4804 54596 4856 54602
rect 4804 54538 4856 54544
rect 4816 54330 4844 54538
rect 4804 54324 4856 54330
rect 4804 54266 4856 54272
rect 4988 53440 5040 53446
rect 4988 53382 5040 53388
rect 5000 53242 5028 53382
rect 4988 53236 5040 53242
rect 4988 53178 5040 53184
rect 4436 53032 4488 53038
rect 4436 52974 4488 52980
rect 2350 52796 2658 52805
rect 2350 52794 2356 52796
rect 2412 52794 2436 52796
rect 2492 52794 2516 52796
rect 2572 52794 2596 52796
rect 2652 52794 2658 52796
rect 2412 52742 2414 52794
rect 2594 52742 2596 52794
rect 2350 52740 2356 52742
rect 2412 52740 2436 52742
rect 2492 52740 2516 52742
rect 2572 52740 2596 52742
rect 2652 52740 2658 52742
rect 2350 52731 2658 52740
rect 3010 52252 3318 52261
rect 3010 52250 3016 52252
rect 3072 52250 3096 52252
rect 3152 52250 3176 52252
rect 3232 52250 3256 52252
rect 3312 52250 3318 52252
rect 3072 52198 3074 52250
rect 3254 52198 3256 52250
rect 3010 52196 3016 52198
rect 3072 52196 3096 52198
rect 3152 52196 3176 52198
rect 3232 52196 3256 52198
rect 3312 52196 3318 52198
rect 3010 52187 3318 52196
rect 4448 51950 4476 52974
rect 4436 51944 4488 51950
rect 4436 51886 4488 51892
rect 4712 51944 4764 51950
rect 4712 51886 4764 51892
rect 2350 51708 2658 51717
rect 2350 51706 2356 51708
rect 2412 51706 2436 51708
rect 2492 51706 2516 51708
rect 2572 51706 2596 51708
rect 2652 51706 2658 51708
rect 2412 51654 2414 51706
rect 2594 51654 2596 51706
rect 2350 51652 2356 51654
rect 2412 51652 2436 51654
rect 2492 51652 2516 51654
rect 2572 51652 2596 51654
rect 2652 51652 2658 51654
rect 2350 51643 2658 51652
rect 3010 51164 3318 51173
rect 3010 51162 3016 51164
rect 3072 51162 3096 51164
rect 3152 51162 3176 51164
rect 3232 51162 3256 51164
rect 3312 51162 3318 51164
rect 3072 51110 3074 51162
rect 3254 51110 3256 51162
rect 3010 51108 3016 51110
rect 3072 51108 3096 51110
rect 3152 51108 3176 51110
rect 3232 51108 3256 51110
rect 3312 51108 3318 51110
rect 3010 51099 3318 51108
rect 2350 50620 2658 50629
rect 2350 50618 2356 50620
rect 2412 50618 2436 50620
rect 2492 50618 2516 50620
rect 2572 50618 2596 50620
rect 2652 50618 2658 50620
rect 2412 50566 2414 50618
rect 2594 50566 2596 50618
rect 2350 50564 2356 50566
rect 2412 50564 2436 50566
rect 2492 50564 2516 50566
rect 2572 50564 2596 50566
rect 2652 50564 2658 50566
rect 2350 50555 2658 50564
rect 4448 50318 4476 51886
rect 4724 51610 4752 51886
rect 4712 51604 4764 51610
rect 4712 51546 4764 51552
rect 4896 50720 4948 50726
rect 4896 50662 4948 50668
rect 4908 50386 4936 50662
rect 4896 50380 4948 50386
rect 4896 50322 4948 50328
rect 4436 50312 4488 50318
rect 4436 50254 4488 50260
rect 3010 50076 3318 50085
rect 3010 50074 3016 50076
rect 3072 50074 3096 50076
rect 3152 50074 3176 50076
rect 3232 50074 3256 50076
rect 3312 50074 3318 50076
rect 3072 50022 3074 50074
rect 3254 50022 3256 50074
rect 3010 50020 3016 50022
rect 3072 50020 3096 50022
rect 3152 50020 3176 50022
rect 3232 50020 3256 50022
rect 3312 50020 3318 50022
rect 3010 50011 3318 50020
rect 4448 49774 4476 50254
rect 5552 49842 5580 65010
rect 5828 63918 5856 65554
rect 6104 65550 6132 66574
rect 6092 65544 6144 65550
rect 6092 65486 6144 65492
rect 5908 63980 5960 63986
rect 5908 63922 5960 63928
rect 5724 63912 5776 63918
rect 5724 63854 5776 63860
rect 5816 63912 5868 63918
rect 5816 63854 5868 63860
rect 5736 63578 5764 63854
rect 5724 63572 5776 63578
rect 5724 63514 5776 63520
rect 5736 63034 5764 63514
rect 5828 63186 5856 63854
rect 5920 63306 5948 63922
rect 5908 63300 5960 63306
rect 5908 63242 5960 63248
rect 5828 63158 5948 63186
rect 5724 63028 5776 63034
rect 5724 62970 5776 62976
rect 5920 62830 5948 63158
rect 5908 62824 5960 62830
rect 5908 62766 5960 62772
rect 6092 62824 6144 62830
rect 6092 62766 6144 62772
rect 5724 61056 5776 61062
rect 5724 60998 5776 61004
rect 5736 60734 5764 60998
rect 5644 60722 5764 60734
rect 5632 60716 5764 60722
rect 5684 60706 5764 60716
rect 5632 60658 5684 60664
rect 5736 60042 5764 60706
rect 5920 60654 5948 62766
rect 6104 62150 6132 62766
rect 6092 62144 6144 62150
rect 6092 62086 6144 62092
rect 6104 61878 6132 62086
rect 6092 61872 6144 61878
rect 6092 61814 6144 61820
rect 6104 60858 6132 61814
rect 6092 60852 6144 60858
rect 6092 60794 6144 60800
rect 5908 60648 5960 60654
rect 5908 60590 5960 60596
rect 5920 60178 5948 60590
rect 5908 60172 5960 60178
rect 5908 60114 5960 60120
rect 5724 60036 5776 60042
rect 5724 59978 5776 59984
rect 5724 59424 5776 59430
rect 5724 59366 5776 59372
rect 5736 58546 5764 59366
rect 5920 59090 5948 60114
rect 6184 59968 6236 59974
rect 6184 59910 6236 59916
rect 6196 59430 6224 59910
rect 6184 59424 6236 59430
rect 6184 59366 6236 59372
rect 6196 59090 6224 59366
rect 5908 59084 5960 59090
rect 5908 59026 5960 59032
rect 6184 59084 6236 59090
rect 6184 59026 6236 59032
rect 5724 58540 5776 58546
rect 5724 58482 5776 58488
rect 5736 57526 5764 58482
rect 5724 57520 5776 57526
rect 5724 57462 5776 57468
rect 5920 56914 5948 59026
rect 6000 58880 6052 58886
rect 6000 58822 6052 58828
rect 6012 58342 6040 58822
rect 6000 58336 6052 58342
rect 6000 58278 6052 58284
rect 6012 57798 6040 58278
rect 6000 57792 6052 57798
rect 6000 57734 6052 57740
rect 5908 56908 5960 56914
rect 5908 56850 5960 56856
rect 5632 56704 5684 56710
rect 5632 56646 5684 56652
rect 5644 56438 5672 56646
rect 5632 56432 5684 56438
rect 5632 56374 5684 56380
rect 5920 56302 5948 56850
rect 6012 56846 6040 57734
rect 6092 57248 6144 57254
rect 6092 57190 6144 57196
rect 6184 57248 6236 57254
rect 6184 57190 6236 57196
rect 6104 56914 6132 57190
rect 6092 56908 6144 56914
rect 6092 56850 6144 56856
rect 6000 56840 6052 56846
rect 6000 56782 6052 56788
rect 6196 56438 6224 57190
rect 6288 57050 6316 68818
rect 6368 67040 6420 67046
rect 6368 66982 6420 66988
rect 6380 66298 6408 66982
rect 6368 66292 6420 66298
rect 6368 66234 6420 66240
rect 6472 65498 6500 70366
rect 6564 70366 6684 70394
rect 6564 68490 6592 70366
rect 6644 69216 6696 69222
rect 6644 69158 6696 69164
rect 6656 68814 6684 69158
rect 6748 68814 6776 70450
rect 6932 70106 6960 70926
rect 7012 70848 7064 70854
rect 7012 70790 7064 70796
rect 7024 70582 7052 70790
rect 7116 70582 7144 71946
rect 7012 70576 7064 70582
rect 7012 70518 7064 70524
rect 7104 70576 7156 70582
rect 7104 70518 7156 70524
rect 7012 70440 7064 70446
rect 7012 70382 7064 70388
rect 6920 70100 6972 70106
rect 6920 70042 6972 70048
rect 6644 68808 6696 68814
rect 6644 68750 6696 68756
rect 6736 68808 6788 68814
rect 6736 68750 6788 68756
rect 6564 68462 6684 68490
rect 6552 68332 6604 68338
rect 6552 68274 6604 68280
rect 6564 67930 6592 68274
rect 6552 67924 6604 67930
rect 6552 67866 6604 67872
rect 6564 67386 6592 67866
rect 6552 67380 6604 67386
rect 6552 67322 6604 67328
rect 6656 65498 6684 68462
rect 6748 67726 6776 68750
rect 6828 68264 6880 68270
rect 6828 68206 6880 68212
rect 6736 67720 6788 67726
rect 6736 67662 6788 67668
rect 6748 66570 6776 67662
rect 6840 67182 6868 68206
rect 7024 67794 7052 70382
rect 7116 69426 7144 70518
rect 7104 69420 7156 69426
rect 7104 69362 7156 69368
rect 7116 68746 7144 69362
rect 7104 68740 7156 68746
rect 7104 68682 7156 68688
rect 7012 67788 7064 67794
rect 7012 67730 7064 67736
rect 7116 67658 7144 68682
rect 7012 67652 7064 67658
rect 7012 67594 7064 67600
rect 7104 67652 7156 67658
rect 7104 67594 7156 67600
rect 7024 67386 7052 67594
rect 7012 67380 7064 67386
rect 7012 67322 7064 67328
rect 6920 67312 6972 67318
rect 6920 67254 6972 67260
rect 6828 67176 6880 67182
rect 6828 67118 6880 67124
rect 6736 66564 6788 66570
rect 6736 66506 6788 66512
rect 6748 66094 6776 66506
rect 6736 66088 6788 66094
rect 6736 66030 6788 66036
rect 6380 65470 6500 65498
rect 6564 65470 6684 65498
rect 6276 57044 6328 57050
rect 6276 56986 6328 56992
rect 6288 56846 6316 56986
rect 6276 56840 6328 56846
rect 6276 56782 6328 56788
rect 6184 56432 6236 56438
rect 6184 56374 6236 56380
rect 5632 56296 5684 56302
rect 5632 56238 5684 56244
rect 5908 56296 5960 56302
rect 5908 56238 5960 56244
rect 5644 55622 5672 56238
rect 5908 55752 5960 55758
rect 6288 55706 6316 56782
rect 6380 56370 6408 65470
rect 6460 64456 6512 64462
rect 6460 64398 6512 64404
rect 6472 63578 6500 64398
rect 6460 63572 6512 63578
rect 6460 63514 6512 63520
rect 6460 62280 6512 62286
rect 6460 62222 6512 62228
rect 6472 61946 6500 62222
rect 6460 61940 6512 61946
rect 6460 61882 6512 61888
rect 6460 59628 6512 59634
rect 6460 59570 6512 59576
rect 6472 59226 6500 59570
rect 6460 59220 6512 59226
rect 6460 59162 6512 59168
rect 6460 58540 6512 58546
rect 6460 58482 6512 58488
rect 6472 58138 6500 58482
rect 6460 58132 6512 58138
rect 6460 58074 6512 58080
rect 6460 57860 6512 57866
rect 6460 57802 6512 57808
rect 6472 56506 6500 57802
rect 6460 56500 6512 56506
rect 6460 56442 6512 56448
rect 6368 56364 6420 56370
rect 6368 56306 6420 56312
rect 5908 55694 5960 55700
rect 5632 55616 5684 55622
rect 5632 55558 5684 55564
rect 5644 54330 5672 55558
rect 5920 54670 5948 55694
rect 6196 55678 6316 55706
rect 5908 54664 5960 54670
rect 5908 54606 5960 54612
rect 5816 54528 5868 54534
rect 5816 54470 5868 54476
rect 5632 54324 5684 54330
rect 5632 54266 5684 54272
rect 5828 53990 5856 54470
rect 5816 53984 5868 53990
rect 5816 53926 5868 53932
rect 5828 53514 5856 53926
rect 5816 53508 5868 53514
rect 5816 53450 5868 53456
rect 5920 53038 5948 54606
rect 6196 54126 6224 55678
rect 6276 55616 6328 55622
rect 6276 55558 6328 55564
rect 6288 55418 6316 55558
rect 6276 55412 6328 55418
rect 6276 55354 6328 55360
rect 6276 55276 6328 55282
rect 6276 55218 6328 55224
rect 6184 54120 6236 54126
rect 6184 54062 6236 54068
rect 6196 53650 6224 54062
rect 6184 53644 6236 53650
rect 6184 53586 6236 53592
rect 6184 53440 6236 53446
rect 6184 53382 6236 53388
rect 5908 53032 5960 53038
rect 5960 52980 6132 52986
rect 5908 52974 6132 52980
rect 5920 52958 6132 52974
rect 5724 51808 5776 51814
rect 5724 51750 5776 51756
rect 5736 51474 5764 51750
rect 5724 51468 5776 51474
rect 5724 51410 5776 51416
rect 5908 51468 5960 51474
rect 5908 51410 5960 51416
rect 5736 50930 5764 51410
rect 5724 50924 5776 50930
rect 5724 50866 5776 50872
rect 5920 50862 5948 51410
rect 5816 50856 5868 50862
rect 5816 50798 5868 50804
rect 5908 50856 5960 50862
rect 5908 50798 5960 50804
rect 5724 50720 5776 50726
rect 5724 50662 5776 50668
rect 5540 49836 5592 49842
rect 5540 49778 5592 49784
rect 4436 49768 4488 49774
rect 4436 49710 4488 49716
rect 2350 49532 2658 49541
rect 2350 49530 2356 49532
rect 2412 49530 2436 49532
rect 2492 49530 2516 49532
rect 2572 49530 2596 49532
rect 2652 49530 2658 49532
rect 2412 49478 2414 49530
rect 2594 49478 2596 49530
rect 2350 49476 2356 49478
rect 2412 49476 2436 49478
rect 2492 49476 2516 49478
rect 2572 49476 2596 49478
rect 2652 49476 2658 49478
rect 2350 49467 2658 49476
rect 4448 49230 4476 49710
rect 4436 49224 4488 49230
rect 4436 49166 4488 49172
rect 3010 48988 3318 48997
rect 3010 48986 3016 48988
rect 3072 48986 3096 48988
rect 3152 48986 3176 48988
rect 3232 48986 3256 48988
rect 3312 48986 3318 48988
rect 3072 48934 3074 48986
rect 3254 48934 3256 48986
rect 3010 48932 3016 48934
rect 3072 48932 3096 48934
rect 3152 48932 3176 48934
rect 3232 48932 3256 48934
rect 3312 48932 3318 48934
rect 3010 48923 3318 48932
rect 2350 48444 2658 48453
rect 2350 48442 2356 48444
rect 2412 48442 2436 48444
rect 2492 48442 2516 48444
rect 2572 48442 2596 48444
rect 2652 48442 2658 48444
rect 2412 48390 2414 48442
rect 2594 48390 2596 48442
rect 2350 48388 2356 48390
rect 2412 48388 2436 48390
rect 2492 48388 2516 48390
rect 2572 48388 2596 48390
rect 2652 48388 2658 48390
rect 2350 48379 2658 48388
rect 3010 47900 3318 47909
rect 3010 47898 3016 47900
rect 3072 47898 3096 47900
rect 3152 47898 3176 47900
rect 3232 47898 3256 47900
rect 3312 47898 3318 47900
rect 3072 47846 3074 47898
rect 3254 47846 3256 47898
rect 3010 47844 3016 47846
rect 3072 47844 3096 47846
rect 3152 47844 3176 47846
rect 3232 47844 3256 47846
rect 3312 47844 3318 47846
rect 3010 47835 3318 47844
rect 4448 47598 4476 49166
rect 4988 49156 5040 49162
rect 4988 49098 5040 49104
rect 5000 48890 5028 49098
rect 4988 48884 5040 48890
rect 4988 48826 5040 48832
rect 4896 48000 4948 48006
rect 4896 47942 4948 47948
rect 4908 47802 4936 47942
rect 4896 47796 4948 47802
rect 4896 47738 4948 47744
rect 4436 47592 4488 47598
rect 4436 47534 4488 47540
rect 2350 47356 2658 47365
rect 2350 47354 2356 47356
rect 2412 47354 2436 47356
rect 2492 47354 2516 47356
rect 2572 47354 2596 47356
rect 2652 47354 2658 47356
rect 2412 47302 2414 47354
rect 2594 47302 2596 47354
rect 2350 47300 2356 47302
rect 2412 47300 2436 47302
rect 2492 47300 2516 47302
rect 2572 47300 2596 47302
rect 2652 47300 2658 47302
rect 2350 47291 2658 47300
rect 3010 46812 3318 46821
rect 3010 46810 3016 46812
rect 3072 46810 3096 46812
rect 3152 46810 3176 46812
rect 3232 46810 3256 46812
rect 3312 46810 3318 46812
rect 3072 46758 3074 46810
rect 3254 46758 3256 46810
rect 3010 46756 3016 46758
rect 3072 46756 3096 46758
rect 3152 46756 3176 46758
rect 3232 46756 3256 46758
rect 3312 46756 3318 46758
rect 3010 46747 3318 46756
rect 4448 46510 4476 47534
rect 5448 46912 5500 46918
rect 5448 46854 5500 46860
rect 4436 46504 4488 46510
rect 4436 46446 4488 46452
rect 4712 46504 4764 46510
rect 4712 46446 4764 46452
rect 2350 46268 2658 46277
rect 2350 46266 2356 46268
rect 2412 46266 2436 46268
rect 2492 46266 2516 46268
rect 2572 46266 2596 46268
rect 2652 46266 2658 46268
rect 2412 46214 2414 46266
rect 2594 46214 2596 46266
rect 2350 46212 2356 46214
rect 2412 46212 2436 46214
rect 2492 46212 2516 46214
rect 2572 46212 2596 46214
rect 2652 46212 2658 46214
rect 2350 46203 2658 46212
rect 3010 45724 3318 45733
rect 3010 45722 3016 45724
rect 3072 45722 3096 45724
rect 3152 45722 3176 45724
rect 3232 45722 3256 45724
rect 3312 45722 3318 45724
rect 3072 45670 3074 45722
rect 3254 45670 3256 45722
rect 3010 45668 3016 45670
rect 3072 45668 3096 45670
rect 3152 45668 3176 45670
rect 3232 45668 3256 45670
rect 3312 45668 3318 45670
rect 3010 45659 3318 45668
rect 4448 45286 4476 46446
rect 4724 46170 4752 46446
rect 4712 46164 4764 46170
rect 4712 46106 4764 46112
rect 5460 45966 5488 46854
rect 5448 45960 5500 45966
rect 5448 45902 5500 45908
rect 4620 45416 4672 45422
rect 4620 45358 4672 45364
rect 4436 45280 4488 45286
rect 4436 45222 4488 45228
rect 2350 45180 2658 45189
rect 2350 45178 2356 45180
rect 2412 45178 2436 45180
rect 2492 45178 2516 45180
rect 2572 45178 2596 45180
rect 2652 45178 2658 45180
rect 2412 45126 2414 45178
rect 2594 45126 2596 45178
rect 2350 45124 2356 45126
rect 2412 45124 2436 45126
rect 2492 45124 2516 45126
rect 2572 45124 2596 45126
rect 2652 45124 2658 45126
rect 2350 45115 2658 45124
rect 3010 44636 3318 44645
rect 3010 44634 3016 44636
rect 3072 44634 3096 44636
rect 3152 44634 3176 44636
rect 3232 44634 3256 44636
rect 3312 44634 3318 44636
rect 3072 44582 3074 44634
rect 3254 44582 3256 44634
rect 3010 44580 3016 44582
rect 3072 44580 3096 44582
rect 3152 44580 3176 44582
rect 3232 44580 3256 44582
rect 3312 44580 3318 44582
rect 3010 44571 3318 44580
rect 2350 44092 2658 44101
rect 2350 44090 2356 44092
rect 2412 44090 2436 44092
rect 2492 44090 2516 44092
rect 2572 44090 2596 44092
rect 2652 44090 2658 44092
rect 2412 44038 2414 44090
rect 2594 44038 2596 44090
rect 2350 44036 2356 44038
rect 2412 44036 2436 44038
rect 2492 44036 2516 44038
rect 2572 44036 2596 44038
rect 2652 44036 2658 44038
rect 2350 44027 2658 44036
rect 4448 43790 4476 45222
rect 4632 45082 4660 45358
rect 4620 45076 4672 45082
rect 4620 45018 4672 45024
rect 5356 44396 5408 44402
rect 5356 44338 5408 44344
rect 5172 44192 5224 44198
rect 5172 44134 5224 44140
rect 5184 43858 5212 44134
rect 5172 43852 5224 43858
rect 5172 43794 5224 43800
rect 4436 43784 4488 43790
rect 4436 43726 4488 43732
rect 3010 43548 3318 43557
rect 3010 43546 3016 43548
rect 3072 43546 3096 43548
rect 3152 43546 3176 43548
rect 3232 43546 3256 43548
rect 3312 43546 3318 43548
rect 3072 43494 3074 43546
rect 3254 43494 3256 43546
rect 3010 43492 3016 43494
rect 3072 43492 3096 43494
rect 3152 43492 3176 43494
rect 3232 43492 3256 43494
rect 3312 43492 3318 43494
rect 3010 43483 3318 43492
rect 2350 43004 2658 43013
rect 2350 43002 2356 43004
rect 2412 43002 2436 43004
rect 2492 43002 2516 43004
rect 2572 43002 2596 43004
rect 2652 43002 2658 43004
rect 2412 42950 2414 43002
rect 2594 42950 2596 43002
rect 2350 42948 2356 42950
rect 2412 42948 2436 42950
rect 2492 42948 2516 42950
rect 2572 42948 2596 42950
rect 2652 42948 2658 42950
rect 2350 42939 2658 42948
rect 4448 42702 4476 43726
rect 5368 43450 5396 44338
rect 5356 43444 5408 43450
rect 5356 43386 5408 43392
rect 4436 42696 4488 42702
rect 4436 42638 4488 42644
rect 3010 42460 3318 42469
rect 3010 42458 3016 42460
rect 3072 42458 3096 42460
rect 3152 42458 3176 42460
rect 3232 42458 3256 42460
rect 3312 42458 3318 42460
rect 3072 42406 3074 42458
rect 3254 42406 3256 42458
rect 3010 42404 3016 42406
rect 3072 42404 3096 42406
rect 3152 42404 3176 42406
rect 3232 42404 3256 42406
rect 3312 42404 3318 42406
rect 3010 42395 3318 42404
rect 2350 41916 2658 41925
rect 2350 41914 2356 41916
rect 2412 41914 2436 41916
rect 2492 41914 2516 41916
rect 2572 41914 2596 41916
rect 2652 41914 2658 41916
rect 2412 41862 2414 41914
rect 2594 41862 2596 41914
rect 2350 41860 2356 41862
rect 2412 41860 2436 41862
rect 2492 41860 2516 41862
rect 2572 41860 2596 41862
rect 2652 41860 2658 41862
rect 2350 41851 2658 41860
rect 3010 41372 3318 41381
rect 3010 41370 3016 41372
rect 3072 41370 3096 41372
rect 3152 41370 3176 41372
rect 3232 41370 3256 41372
rect 3312 41370 3318 41372
rect 3072 41318 3074 41370
rect 3254 41318 3256 41370
rect 3010 41316 3016 41318
rect 3072 41316 3096 41318
rect 3152 41316 3176 41318
rect 3232 41316 3256 41318
rect 3312 41316 3318 41318
rect 3010 41307 3318 41316
rect 4448 41138 4476 42638
rect 4988 42628 5040 42634
rect 4988 42570 5040 42576
rect 5000 42362 5028 42570
rect 4988 42356 5040 42362
rect 4988 42298 5040 42304
rect 4436 41132 4488 41138
rect 4436 41074 4488 41080
rect 4712 41064 4764 41070
rect 4712 41006 4764 41012
rect 2350 40828 2658 40837
rect 2350 40826 2356 40828
rect 2412 40826 2436 40828
rect 2492 40826 2516 40828
rect 2572 40826 2596 40828
rect 2652 40826 2658 40828
rect 2412 40774 2414 40826
rect 2594 40774 2596 40826
rect 2350 40772 2356 40774
rect 2412 40772 2436 40774
rect 2492 40772 2516 40774
rect 2572 40772 2596 40774
rect 2652 40772 2658 40774
rect 2350 40763 2658 40772
rect 4724 40730 4752 41006
rect 4712 40724 4764 40730
rect 4712 40666 4764 40672
rect 4804 40520 4856 40526
rect 4804 40462 4856 40468
rect 3010 40284 3318 40293
rect 3010 40282 3016 40284
rect 3072 40282 3096 40284
rect 3152 40282 3176 40284
rect 3232 40282 3256 40284
rect 3312 40282 3318 40284
rect 3072 40230 3074 40282
rect 3254 40230 3256 40282
rect 3010 40228 3016 40230
rect 3072 40228 3096 40230
rect 3152 40228 3176 40230
rect 3232 40228 3256 40230
rect 3312 40228 3318 40230
rect 3010 40219 3318 40228
rect 4816 40186 4844 40462
rect 5552 40390 5580 49778
rect 5736 45830 5764 50662
rect 5828 50522 5856 50798
rect 5816 50516 5868 50522
rect 5816 50458 5868 50464
rect 5828 48890 5856 50458
rect 5920 49178 5948 50798
rect 5920 49150 6040 49178
rect 5908 49088 5960 49094
rect 5908 49030 5960 49036
rect 5816 48884 5868 48890
rect 5816 48826 5868 48832
rect 5920 48686 5948 49030
rect 6012 48686 6040 49150
rect 5908 48680 5960 48686
rect 5908 48622 5960 48628
rect 6000 48680 6052 48686
rect 6000 48622 6052 48628
rect 5920 48142 5948 48622
rect 6012 48210 6040 48622
rect 6000 48204 6052 48210
rect 6000 48146 6052 48152
rect 5908 48136 5960 48142
rect 5908 48078 5960 48084
rect 6012 47122 6040 48146
rect 6104 47734 6132 52958
rect 6196 52902 6224 53382
rect 6184 52896 6236 52902
rect 6184 52838 6236 52844
rect 6196 52494 6224 52838
rect 6184 52488 6236 52494
rect 6184 52430 6236 52436
rect 6196 51406 6224 52430
rect 6184 51400 6236 51406
rect 6184 51342 6236 51348
rect 6184 48000 6236 48006
rect 6184 47942 6236 47948
rect 6092 47728 6144 47734
rect 6092 47670 6144 47676
rect 6000 47116 6052 47122
rect 6000 47058 6052 47064
rect 6012 46034 6040 47058
rect 6104 46986 6132 47670
rect 6196 47462 6224 47942
rect 6184 47456 6236 47462
rect 6184 47398 6236 47404
rect 6196 47122 6224 47398
rect 6184 47116 6236 47122
rect 6184 47058 6236 47064
rect 6092 46980 6144 46986
rect 6092 46922 6144 46928
rect 6184 46912 6236 46918
rect 6184 46854 6236 46860
rect 6196 46510 6224 46854
rect 6184 46504 6236 46510
rect 6184 46446 6236 46452
rect 6000 46028 6052 46034
rect 6000 45970 6052 45976
rect 5632 45824 5684 45830
rect 5632 45766 5684 45772
rect 5724 45824 5776 45830
rect 5724 45766 5776 45772
rect 5644 44878 5672 45766
rect 5632 44872 5684 44878
rect 5632 44814 5684 44820
rect 6012 43246 6040 45970
rect 6196 45966 6224 46446
rect 6184 45960 6236 45966
rect 6184 45902 6236 45908
rect 6092 45824 6144 45830
rect 6092 45766 6144 45772
rect 6104 45626 6132 45766
rect 6092 45620 6144 45626
rect 6092 45562 6144 45568
rect 6288 43994 6316 55218
rect 6276 43988 6328 43994
rect 6276 43930 6328 43936
rect 6288 43450 6316 43930
rect 6276 43444 6328 43450
rect 6276 43386 6328 43392
rect 6184 43308 6236 43314
rect 6184 43250 6236 43256
rect 6000 43240 6052 43246
rect 6000 43182 6052 43188
rect 6012 42378 6040 43182
rect 5920 42350 6040 42378
rect 5920 42294 5948 42350
rect 6196 42294 6224 43250
rect 5908 42288 5960 42294
rect 6184 42288 6236 42294
rect 5908 42230 5960 42236
rect 6104 42236 6184 42242
rect 6104 42230 6236 42236
rect 5920 41818 5948 42230
rect 6104 42214 6224 42230
rect 5908 41812 5960 41818
rect 5908 41754 5960 41760
rect 5540 40384 5592 40390
rect 5540 40326 5592 40332
rect 4804 40180 4856 40186
rect 4804 40122 4856 40128
rect 5632 40112 5684 40118
rect 5630 40080 5632 40089
rect 5684 40080 5686 40089
rect 5630 40015 5686 40024
rect 5920 39982 5948 41754
rect 6104 41274 6132 42214
rect 6184 41540 6236 41546
rect 6184 41482 6236 41488
rect 6196 41449 6224 41482
rect 6182 41440 6238 41449
rect 6182 41375 6238 41384
rect 6092 41268 6144 41274
rect 6092 41210 6144 41216
rect 6104 40186 6132 41210
rect 6380 40186 6408 56306
rect 6472 55894 6500 56442
rect 6460 55888 6512 55894
rect 6460 55830 6512 55836
rect 6460 55752 6512 55758
rect 6460 55694 6512 55700
rect 6472 55418 6500 55694
rect 6460 55412 6512 55418
rect 6460 55354 6512 55360
rect 6460 54188 6512 54194
rect 6460 54130 6512 54136
rect 6472 53786 6500 54130
rect 6460 53780 6512 53786
rect 6460 53722 6512 53728
rect 6460 53100 6512 53106
rect 6460 53042 6512 53048
rect 6472 52698 6500 53042
rect 6460 52692 6512 52698
rect 6460 52634 6512 52640
rect 6460 51400 6512 51406
rect 6460 51342 6512 51348
rect 6472 51066 6500 51342
rect 6460 51060 6512 51066
rect 6460 51002 6512 51008
rect 6564 50726 6592 65470
rect 6748 64462 6776 66030
rect 6840 65618 6868 67118
rect 6932 66842 6960 67254
rect 6920 66836 6972 66842
rect 6920 66778 6972 66784
rect 6828 65612 6880 65618
rect 6828 65554 6880 65560
rect 6932 65550 6960 66778
rect 7012 66632 7064 66638
rect 7012 66574 7064 66580
rect 7104 66632 7156 66638
rect 7104 66574 7156 66580
rect 7024 66230 7052 66574
rect 7012 66224 7064 66230
rect 7012 66166 7064 66172
rect 7116 66042 7144 66574
rect 7024 66014 7144 66042
rect 6920 65544 6972 65550
rect 6920 65486 6972 65492
rect 6920 65408 6972 65414
rect 6920 65350 6972 65356
rect 6932 65210 6960 65350
rect 6920 65204 6972 65210
rect 6920 65146 6972 65152
rect 7024 65090 7052 66014
rect 6932 65062 7052 65090
rect 7104 65068 7156 65074
rect 6736 64456 6788 64462
rect 6736 64398 6788 64404
rect 6644 64320 6696 64326
rect 6644 64262 6696 64268
rect 6656 64122 6684 64262
rect 6644 64116 6696 64122
rect 6644 64058 6696 64064
rect 6748 63782 6776 64398
rect 6736 63776 6788 63782
rect 6736 63718 6788 63724
rect 6644 63232 6696 63238
rect 6644 63174 6696 63180
rect 6656 55282 6684 63174
rect 6748 62286 6776 63718
rect 6736 62280 6788 62286
rect 6736 62222 6788 62228
rect 6748 60654 6776 62222
rect 6932 61305 6960 65062
rect 7104 65010 7156 65016
rect 7012 64864 7064 64870
rect 7012 64806 7064 64812
rect 7024 64530 7052 64806
rect 7012 64524 7064 64530
rect 7012 64466 7064 64472
rect 7012 64116 7064 64122
rect 7012 64058 7064 64064
rect 7024 62354 7052 64058
rect 7116 63510 7144 65010
rect 7104 63504 7156 63510
rect 7104 63446 7156 63452
rect 7104 63300 7156 63306
rect 7104 63242 7156 63248
rect 7116 62490 7144 63242
rect 7104 62484 7156 62490
rect 7104 62426 7156 62432
rect 7012 62348 7064 62354
rect 7012 62290 7064 62296
rect 6918 61296 6974 61305
rect 6918 61231 6974 61240
rect 6828 61192 6880 61198
rect 7024 61146 7052 62290
rect 7104 62144 7156 62150
rect 7104 62086 7156 62092
rect 7116 61946 7144 62086
rect 7104 61940 7156 61946
rect 7104 61882 7156 61888
rect 7104 61600 7156 61606
rect 7104 61542 7156 61548
rect 6828 61134 6880 61140
rect 6736 60648 6788 60654
rect 6736 60590 6788 60596
rect 6748 59566 6776 60590
rect 6840 60314 6868 61134
rect 6932 61130 7052 61146
rect 6920 61124 7052 61130
rect 6972 61118 7052 61124
rect 6920 61066 6972 61072
rect 6932 60790 6960 61066
rect 7116 61062 7144 61542
rect 7012 61056 7064 61062
rect 7012 60998 7064 61004
rect 7104 61056 7156 61062
rect 7104 60998 7156 61004
rect 7024 60790 7052 60998
rect 7104 60852 7156 60858
rect 7104 60794 7156 60800
rect 6920 60784 6972 60790
rect 6920 60726 6972 60732
rect 7012 60784 7064 60790
rect 7012 60726 7064 60732
rect 7012 60648 7064 60654
rect 6932 60596 7012 60602
rect 6932 60590 7064 60596
rect 6932 60574 7052 60590
rect 6828 60308 6880 60314
rect 6828 60250 6880 60256
rect 6736 59560 6788 59566
rect 6736 59502 6788 59508
rect 6748 58478 6776 59502
rect 6736 58472 6788 58478
rect 6736 58414 6788 58420
rect 6828 57452 6880 57458
rect 6828 57394 6880 57400
rect 6736 56908 6788 56914
rect 6736 56850 6788 56856
rect 6748 55826 6776 56850
rect 6840 56506 6868 57394
rect 6828 56500 6880 56506
rect 6828 56442 6880 56448
rect 6932 56386 6960 60574
rect 7012 60512 7064 60518
rect 7012 60454 7064 60460
rect 7024 60110 7052 60454
rect 7012 60104 7064 60110
rect 7012 60046 7064 60052
rect 7012 59968 7064 59974
rect 7012 59910 7064 59916
rect 7024 59158 7052 59910
rect 7116 59566 7144 60794
rect 7104 59560 7156 59566
rect 7104 59502 7156 59508
rect 7104 59424 7156 59430
rect 7104 59366 7156 59372
rect 7012 59152 7064 59158
rect 7012 59094 7064 59100
rect 7024 58002 7052 59094
rect 7116 59022 7144 59366
rect 7104 59016 7156 59022
rect 7104 58958 7156 58964
rect 7104 58336 7156 58342
rect 7104 58278 7156 58284
rect 7012 57996 7064 58002
rect 7012 57938 7064 57944
rect 7116 57934 7144 58278
rect 7104 57928 7156 57934
rect 7104 57870 7156 57876
rect 7104 57452 7156 57458
rect 7104 57394 7156 57400
rect 7012 57248 7064 57254
rect 7012 57190 7064 57196
rect 7024 56914 7052 57190
rect 7116 56914 7144 57394
rect 7012 56908 7064 56914
rect 7012 56850 7064 56856
rect 7104 56908 7156 56914
rect 7104 56850 7156 56856
rect 7116 56506 7144 56850
rect 7104 56500 7156 56506
rect 7104 56442 7156 56448
rect 6932 56358 7144 56386
rect 6920 56296 6972 56302
rect 6920 56238 6972 56244
rect 6828 56228 6880 56234
rect 6828 56170 6880 56176
rect 6736 55820 6788 55826
rect 6736 55762 6788 55768
rect 6644 55276 6696 55282
rect 6644 55218 6696 55224
rect 6748 54194 6776 55762
rect 6736 54188 6788 54194
rect 6736 54130 6788 54136
rect 6644 53644 6696 53650
rect 6644 53586 6696 53592
rect 6552 50720 6604 50726
rect 6552 50662 6604 50668
rect 6460 50312 6512 50318
rect 6460 50254 6512 50260
rect 6552 50312 6604 50318
rect 6552 50254 6604 50260
rect 6472 49434 6500 50254
rect 6564 49774 6592 50254
rect 6552 49768 6604 49774
rect 6552 49710 6604 49716
rect 6460 49428 6512 49434
rect 6460 49370 6512 49376
rect 6564 48686 6592 49710
rect 6656 49178 6684 53586
rect 6748 53106 6776 54130
rect 6736 53100 6788 53106
rect 6736 53042 6788 53048
rect 6748 51474 6776 53042
rect 6736 51468 6788 51474
rect 6736 51410 6788 51416
rect 6748 50318 6776 51410
rect 6736 50312 6788 50318
rect 6736 50254 6788 50260
rect 6656 49150 6776 49178
rect 6644 49088 6696 49094
rect 6644 49030 6696 49036
rect 6656 48890 6684 49030
rect 6644 48884 6696 48890
rect 6644 48826 6696 48832
rect 6552 48680 6604 48686
rect 6552 48622 6604 48628
rect 6460 47660 6512 47666
rect 6460 47602 6512 47608
rect 6472 47258 6500 47602
rect 6564 47598 6592 48622
rect 6552 47592 6604 47598
rect 6552 47534 6604 47540
rect 6460 47252 6512 47258
rect 6460 47194 6512 47200
rect 6460 47048 6512 47054
rect 6460 46990 6512 46996
rect 6472 46646 6500 46990
rect 6460 46640 6512 46646
rect 6460 46582 6512 46588
rect 6472 45490 6500 46582
rect 6564 45966 6592 47534
rect 6552 45960 6604 45966
rect 6552 45902 6604 45908
rect 6460 45484 6512 45490
rect 6460 45426 6512 45432
rect 6472 43790 6500 45426
rect 6564 44878 6592 45902
rect 6552 44872 6604 44878
rect 6552 44814 6604 44820
rect 6460 43784 6512 43790
rect 6460 43726 6512 43732
rect 6472 42702 6500 43726
rect 6564 42770 6592 44814
rect 6552 42764 6604 42770
rect 6552 42706 6604 42712
rect 6460 42696 6512 42702
rect 6460 42638 6512 42644
rect 6748 41614 6776 49150
rect 6840 48314 6868 56170
rect 6932 55214 6960 56238
rect 6920 55208 6972 55214
rect 6920 55150 6972 55156
rect 6932 53650 6960 55150
rect 7012 53984 7064 53990
rect 7012 53926 7064 53932
rect 6920 53644 6972 53650
rect 6920 53586 6972 53592
rect 6932 52630 6960 53586
rect 7024 53582 7052 53926
rect 7012 53576 7064 53582
rect 7012 53518 7064 53524
rect 6920 52624 6972 52630
rect 6920 52566 6972 52572
rect 6932 50862 6960 52566
rect 7116 51610 7144 56358
rect 7104 51604 7156 51610
rect 7104 51546 7156 51552
rect 7012 51468 7064 51474
rect 7012 51410 7064 51416
rect 6920 50856 6972 50862
rect 6920 50798 6972 50804
rect 7024 50266 7052 51410
rect 7104 50720 7156 50726
rect 7104 50662 7156 50668
rect 6932 50238 7052 50266
rect 6932 50182 6960 50238
rect 6920 50176 6972 50182
rect 6920 50118 6972 50124
rect 7012 49700 7064 49706
rect 7012 49642 7064 49648
rect 7024 49230 7052 49642
rect 7116 49298 7144 50662
rect 7104 49292 7156 49298
rect 7104 49234 7156 49240
rect 7012 49224 7064 49230
rect 7012 49166 7064 49172
rect 7104 48680 7156 48686
rect 7104 48622 7156 48628
rect 6840 48286 6960 48314
rect 6828 46368 6880 46374
rect 6828 46310 6880 46316
rect 6840 46170 6868 46310
rect 6828 46164 6880 46170
rect 6828 46106 6880 46112
rect 6932 45490 6960 48286
rect 7116 48278 7144 48622
rect 7104 48272 7156 48278
rect 7104 48214 7156 48220
rect 7116 47818 7144 48214
rect 7024 47790 7144 47818
rect 7024 47258 7052 47790
rect 7104 47728 7156 47734
rect 7104 47670 7156 47676
rect 7012 47252 7064 47258
rect 7012 47194 7064 47200
rect 7116 47054 7144 47670
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 7208 45642 7236 79206
rect 7392 79098 7420 79206
rect 7470 79200 7526 80000
rect 7484 79098 7512 79200
rect 7392 79070 7512 79098
rect 7350 77820 7658 77829
rect 7350 77818 7356 77820
rect 7412 77818 7436 77820
rect 7492 77818 7516 77820
rect 7572 77818 7596 77820
rect 7652 77818 7658 77820
rect 7412 77766 7414 77818
rect 7594 77766 7596 77818
rect 7350 77764 7356 77766
rect 7412 77764 7436 77766
rect 7492 77764 7516 77766
rect 7572 77764 7596 77766
rect 7652 77764 7658 77766
rect 7350 77755 7658 77764
rect 8010 77276 8318 77285
rect 8010 77274 8016 77276
rect 8072 77274 8096 77276
rect 8152 77274 8176 77276
rect 8232 77274 8256 77276
rect 8312 77274 8318 77276
rect 8072 77222 8074 77274
rect 8254 77222 8256 77274
rect 8010 77220 8016 77222
rect 8072 77220 8096 77222
rect 8152 77220 8176 77222
rect 8232 77220 8256 77222
rect 8312 77220 8318 77222
rect 8010 77211 8318 77220
rect 7350 76732 7658 76741
rect 7350 76730 7356 76732
rect 7412 76730 7436 76732
rect 7492 76730 7516 76732
rect 7572 76730 7596 76732
rect 7652 76730 7658 76732
rect 7412 76678 7414 76730
rect 7594 76678 7596 76730
rect 7350 76676 7356 76678
rect 7412 76676 7436 76678
rect 7492 76676 7516 76678
rect 7572 76676 7596 76678
rect 7652 76676 7658 76678
rect 7350 76667 7658 76676
rect 8010 76188 8318 76197
rect 8010 76186 8016 76188
rect 8072 76186 8096 76188
rect 8152 76186 8176 76188
rect 8232 76186 8256 76188
rect 8312 76186 8318 76188
rect 8072 76134 8074 76186
rect 8254 76134 8256 76186
rect 8010 76132 8016 76134
rect 8072 76132 8096 76134
rect 8152 76132 8176 76134
rect 8232 76132 8256 76134
rect 8312 76132 8318 76134
rect 8010 76123 8318 76132
rect 7350 75644 7658 75653
rect 7350 75642 7356 75644
rect 7412 75642 7436 75644
rect 7492 75642 7516 75644
rect 7572 75642 7596 75644
rect 7652 75642 7658 75644
rect 7412 75590 7414 75642
rect 7594 75590 7596 75642
rect 7350 75588 7356 75590
rect 7412 75588 7436 75590
rect 7492 75588 7516 75590
rect 7572 75588 7596 75590
rect 7652 75588 7658 75590
rect 7350 75579 7658 75588
rect 8010 75100 8318 75109
rect 8010 75098 8016 75100
rect 8072 75098 8096 75100
rect 8152 75098 8176 75100
rect 8232 75098 8256 75100
rect 8312 75098 8318 75100
rect 8072 75046 8074 75098
rect 8254 75046 8256 75098
rect 8010 75044 8016 75046
rect 8072 75044 8096 75046
rect 8152 75044 8176 75046
rect 8232 75044 8256 75046
rect 8312 75044 8318 75046
rect 8010 75035 8318 75044
rect 7350 74556 7658 74565
rect 7350 74554 7356 74556
rect 7412 74554 7436 74556
rect 7492 74554 7516 74556
rect 7572 74554 7596 74556
rect 7652 74554 7658 74556
rect 7412 74502 7414 74554
rect 7594 74502 7596 74554
rect 7350 74500 7356 74502
rect 7412 74500 7436 74502
rect 7492 74500 7516 74502
rect 7572 74500 7596 74502
rect 7652 74500 7658 74502
rect 7350 74491 7658 74500
rect 7932 74248 7984 74254
rect 7932 74190 7984 74196
rect 7748 73840 7800 73846
rect 7748 73782 7800 73788
rect 7944 73794 7972 74190
rect 8392 74112 8444 74118
rect 8392 74054 8444 74060
rect 8010 74012 8318 74021
rect 8010 74010 8016 74012
rect 8072 74010 8096 74012
rect 8152 74010 8176 74012
rect 8232 74010 8256 74012
rect 8312 74010 8318 74012
rect 8072 73958 8074 74010
rect 8254 73958 8256 74010
rect 8010 73956 8016 73958
rect 8072 73956 8096 73958
rect 8152 73956 8176 73958
rect 8232 73956 8256 73958
rect 8312 73956 8318 73958
rect 8010 73947 8318 73956
rect 7350 73468 7658 73477
rect 7350 73466 7356 73468
rect 7412 73466 7436 73468
rect 7492 73466 7516 73468
rect 7572 73466 7596 73468
rect 7652 73466 7658 73468
rect 7412 73414 7414 73466
rect 7594 73414 7596 73466
rect 7350 73412 7356 73414
rect 7412 73412 7436 73414
rect 7492 73412 7516 73414
rect 7572 73412 7596 73414
rect 7652 73412 7658 73414
rect 7350 73403 7658 73412
rect 7760 73030 7788 73782
rect 7944 73766 8064 73794
rect 8036 73574 8064 73766
rect 8024 73568 8076 73574
rect 8024 73510 8076 73516
rect 7840 73296 7892 73302
rect 7840 73238 7892 73244
rect 7748 73024 7800 73030
rect 7748 72966 7800 72972
rect 7350 72380 7658 72389
rect 7350 72378 7356 72380
rect 7412 72378 7436 72380
rect 7492 72378 7516 72380
rect 7572 72378 7596 72380
rect 7652 72378 7658 72380
rect 7412 72326 7414 72378
rect 7594 72326 7596 72378
rect 7350 72324 7356 72326
rect 7412 72324 7436 72326
rect 7492 72324 7516 72326
rect 7572 72324 7596 72326
rect 7652 72324 7658 72326
rect 7350 72315 7658 72324
rect 7760 71942 7788 72966
rect 7748 71936 7800 71942
rect 7748 71878 7800 71884
rect 7852 71534 7880 73238
rect 8036 73234 8064 73510
rect 8404 73273 8432 74054
rect 8390 73264 8446 73273
rect 8024 73228 8076 73234
rect 8390 73199 8446 73208
rect 8024 73170 8076 73176
rect 7944 73098 8064 73114
rect 7944 73092 8076 73098
rect 7944 73086 8024 73092
rect 7944 72826 7972 73086
rect 8024 73034 8076 73040
rect 8010 72924 8318 72933
rect 8010 72922 8016 72924
rect 8072 72922 8096 72924
rect 8152 72922 8176 72924
rect 8232 72922 8256 72924
rect 8312 72922 8318 72924
rect 8072 72870 8074 72922
rect 8254 72870 8256 72922
rect 8010 72868 8016 72870
rect 8072 72868 8096 72870
rect 8152 72868 8176 72870
rect 8232 72868 8256 72870
rect 8312 72868 8318 72870
rect 8010 72859 8318 72868
rect 7932 72820 7984 72826
rect 7932 72762 7984 72768
rect 7932 71936 7984 71942
rect 7932 71878 7984 71884
rect 8482 71904 8538 71913
rect 7944 71670 7972 71878
rect 8010 71836 8318 71845
rect 8482 71839 8538 71848
rect 8010 71834 8016 71836
rect 8072 71834 8096 71836
rect 8152 71834 8176 71836
rect 8232 71834 8256 71836
rect 8312 71834 8318 71836
rect 8072 71782 8074 71834
rect 8254 71782 8256 71834
rect 8010 71780 8016 71782
rect 8072 71780 8096 71782
rect 8152 71780 8176 71782
rect 8232 71780 8256 71782
rect 8312 71780 8318 71782
rect 8010 71771 8318 71780
rect 8496 71738 8524 71839
rect 8484 71732 8536 71738
rect 8484 71674 8536 71680
rect 7932 71664 7984 71670
rect 7932 71606 7984 71612
rect 7840 71528 7892 71534
rect 7840 71470 7892 71476
rect 7350 71292 7658 71301
rect 7350 71290 7356 71292
rect 7412 71290 7436 71292
rect 7492 71290 7516 71292
rect 7572 71290 7596 71292
rect 7652 71290 7658 71292
rect 7412 71238 7414 71290
rect 7594 71238 7596 71290
rect 7350 71236 7356 71238
rect 7412 71236 7436 71238
rect 7492 71236 7516 71238
rect 7572 71236 7596 71238
rect 7652 71236 7658 71238
rect 7350 71227 7658 71236
rect 7350 70204 7658 70213
rect 7350 70202 7356 70204
rect 7412 70202 7436 70204
rect 7492 70202 7516 70204
rect 7572 70202 7596 70204
rect 7652 70202 7658 70204
rect 7412 70150 7414 70202
rect 7594 70150 7596 70202
rect 7350 70148 7356 70150
rect 7412 70148 7436 70150
rect 7492 70148 7516 70150
rect 7572 70148 7596 70150
rect 7652 70148 7658 70150
rect 7350 70139 7658 70148
rect 7852 69970 7880 71470
rect 7932 70984 7984 70990
rect 7932 70926 7984 70932
rect 7944 70394 7972 70926
rect 8392 70848 8444 70854
rect 8392 70790 8444 70796
rect 8010 70748 8318 70757
rect 8010 70746 8016 70748
rect 8072 70746 8096 70748
rect 8152 70746 8176 70748
rect 8232 70746 8256 70748
rect 8312 70746 8318 70748
rect 8072 70694 8074 70746
rect 8254 70694 8256 70746
rect 8010 70692 8016 70694
rect 8072 70692 8096 70694
rect 8152 70692 8176 70694
rect 8232 70692 8256 70694
rect 8312 70692 8318 70694
rect 8010 70683 8318 70692
rect 8404 70553 8432 70790
rect 8390 70544 8446 70553
rect 8390 70479 8446 70488
rect 7944 70378 8064 70394
rect 7944 70372 8076 70378
rect 7944 70366 8024 70372
rect 7840 69964 7892 69970
rect 7840 69906 7892 69912
rect 7852 69358 7880 69906
rect 7944 69902 7972 70366
rect 8024 70314 8076 70320
rect 7932 69896 7984 69902
rect 7932 69838 7984 69844
rect 8010 69660 8318 69669
rect 8010 69658 8016 69660
rect 8072 69658 8096 69660
rect 8152 69658 8176 69660
rect 8232 69658 8256 69660
rect 8312 69658 8318 69660
rect 8072 69606 8074 69658
rect 8254 69606 8256 69658
rect 8010 69604 8016 69606
rect 8072 69604 8096 69606
rect 8152 69604 8176 69606
rect 8232 69604 8256 69606
rect 8312 69604 8318 69606
rect 8010 69595 8318 69604
rect 8484 69420 8536 69426
rect 8484 69362 8536 69368
rect 7840 69352 7892 69358
rect 7840 69294 7892 69300
rect 7350 69116 7658 69125
rect 7350 69114 7356 69116
rect 7412 69114 7436 69116
rect 7492 69114 7516 69116
rect 7572 69114 7596 69116
rect 7652 69114 7658 69116
rect 7412 69062 7414 69114
rect 7594 69062 7596 69114
rect 7350 69060 7356 69062
rect 7412 69060 7436 69062
rect 7492 69060 7516 69062
rect 7572 69060 7596 69062
rect 7652 69060 7658 69062
rect 7350 69051 7658 69060
rect 7852 68270 7880 69294
rect 8392 69216 8444 69222
rect 8390 69184 8392 69193
rect 8444 69184 8446 69193
rect 8390 69119 8446 69128
rect 8496 69018 8524 69362
rect 8484 69012 8536 69018
rect 8484 68954 8536 68960
rect 8010 68572 8318 68581
rect 8010 68570 8016 68572
rect 8072 68570 8096 68572
rect 8152 68570 8176 68572
rect 8232 68570 8256 68572
rect 8312 68570 8318 68572
rect 8072 68518 8074 68570
rect 8254 68518 8256 68570
rect 8010 68516 8016 68518
rect 8072 68516 8096 68518
rect 8152 68516 8176 68518
rect 8232 68516 8256 68518
rect 8312 68516 8318 68518
rect 8010 68507 8318 68516
rect 7840 68264 7892 68270
rect 7840 68206 7892 68212
rect 7748 68128 7800 68134
rect 7748 68070 7800 68076
rect 7350 68028 7658 68037
rect 7350 68026 7356 68028
rect 7412 68026 7436 68028
rect 7492 68026 7516 68028
rect 7572 68026 7596 68028
rect 7652 68026 7658 68028
rect 7412 67974 7414 68026
rect 7594 67974 7596 68026
rect 7350 67972 7356 67974
rect 7412 67972 7436 67974
rect 7492 67972 7516 67974
rect 7572 67972 7596 67974
rect 7652 67972 7658 67974
rect 7350 67963 7658 67972
rect 7656 67788 7708 67794
rect 7656 67730 7708 67736
rect 7668 67130 7696 67730
rect 7760 67386 7788 68070
rect 7748 67380 7800 67386
rect 7748 67322 7800 67328
rect 7668 67102 7788 67130
rect 7350 66940 7658 66949
rect 7350 66938 7356 66940
rect 7412 66938 7436 66940
rect 7492 66938 7516 66940
rect 7572 66938 7596 66940
rect 7652 66938 7658 66940
rect 7412 66886 7414 66938
rect 7594 66886 7596 66938
rect 7350 66884 7356 66886
rect 7412 66884 7436 66886
rect 7492 66884 7516 66886
rect 7572 66884 7596 66886
rect 7652 66884 7658 66886
rect 7350 66875 7658 66884
rect 7656 66496 7708 66502
rect 7656 66438 7708 66444
rect 7668 66298 7696 66438
rect 7656 66292 7708 66298
rect 7656 66234 7708 66240
rect 7350 65852 7658 65861
rect 7350 65850 7356 65852
rect 7412 65850 7436 65852
rect 7492 65850 7516 65852
rect 7572 65850 7596 65852
rect 7652 65850 7658 65852
rect 7412 65798 7414 65850
rect 7594 65798 7596 65850
rect 7350 65796 7356 65798
rect 7412 65796 7436 65798
rect 7492 65796 7516 65798
rect 7572 65796 7596 65798
rect 7652 65796 7658 65798
rect 7350 65787 7658 65796
rect 7760 65498 7788 67102
rect 7852 66638 7880 68206
rect 8392 68128 8444 68134
rect 8392 68070 8444 68076
rect 8404 67833 8432 68070
rect 8390 67824 8446 67833
rect 8390 67759 8446 67768
rect 8010 67484 8318 67493
rect 8010 67482 8016 67484
rect 8072 67482 8096 67484
rect 8152 67482 8176 67484
rect 8232 67482 8256 67484
rect 8312 67482 8318 67484
rect 8072 67430 8074 67482
rect 8254 67430 8256 67482
rect 8010 67428 8016 67430
rect 8072 67428 8096 67430
rect 8152 67428 8176 67430
rect 8232 67428 8256 67430
rect 8312 67428 8318 67430
rect 8010 67419 8318 67428
rect 8484 67244 8536 67250
rect 8484 67186 8536 67192
rect 8392 67040 8444 67046
rect 8392 66982 8444 66988
rect 7840 66632 7892 66638
rect 7840 66574 7892 66580
rect 8404 66473 8432 66982
rect 8496 66502 8524 67186
rect 8484 66496 8536 66502
rect 8390 66464 8446 66473
rect 8484 66438 8536 66444
rect 8010 66396 8318 66405
rect 8390 66399 8446 66408
rect 8010 66394 8016 66396
rect 8072 66394 8096 66396
rect 8152 66394 8176 66396
rect 8232 66394 8256 66396
rect 8312 66394 8318 66396
rect 8072 66342 8074 66394
rect 8254 66342 8256 66394
rect 8010 66340 8016 66342
rect 8072 66340 8096 66342
rect 8152 66340 8176 66342
rect 8232 66340 8256 66342
rect 8312 66340 8318 66342
rect 8010 66331 8318 66340
rect 8496 66298 8524 66438
rect 8484 66292 8536 66298
rect 8484 66234 8536 66240
rect 7932 65544 7984 65550
rect 7760 65470 7880 65498
rect 7932 65486 7984 65492
rect 7748 65408 7800 65414
rect 7748 65350 7800 65356
rect 7350 64764 7658 64773
rect 7350 64762 7356 64764
rect 7412 64762 7436 64764
rect 7492 64762 7516 64764
rect 7572 64762 7596 64764
rect 7652 64762 7658 64764
rect 7412 64710 7414 64762
rect 7594 64710 7596 64762
rect 7350 64708 7356 64710
rect 7412 64708 7436 64710
rect 7492 64708 7516 64710
rect 7572 64708 7596 64710
rect 7652 64708 7658 64710
rect 7350 64699 7658 64708
rect 7656 64524 7708 64530
rect 7656 64466 7708 64472
rect 7668 64122 7696 64466
rect 7656 64116 7708 64122
rect 7656 64058 7708 64064
rect 7350 63676 7658 63685
rect 7350 63674 7356 63676
rect 7412 63674 7436 63676
rect 7492 63674 7516 63676
rect 7572 63674 7596 63676
rect 7652 63674 7658 63676
rect 7412 63622 7414 63674
rect 7594 63622 7596 63674
rect 7350 63620 7356 63622
rect 7412 63620 7436 63622
rect 7492 63620 7516 63622
rect 7572 63620 7596 63622
rect 7652 63620 7658 63622
rect 7350 63611 7658 63620
rect 7288 63504 7340 63510
rect 7288 63446 7340 63452
rect 7300 63306 7328 63446
rect 7288 63300 7340 63306
rect 7288 63242 7340 63248
rect 7350 62588 7658 62597
rect 7350 62586 7356 62588
rect 7412 62586 7436 62588
rect 7492 62586 7516 62588
rect 7572 62586 7596 62588
rect 7652 62586 7658 62588
rect 7412 62534 7414 62586
rect 7594 62534 7596 62586
rect 7350 62532 7356 62534
rect 7412 62532 7436 62534
rect 7492 62532 7516 62534
rect 7572 62532 7596 62534
rect 7652 62532 7658 62534
rect 7350 62523 7658 62532
rect 7350 61500 7658 61509
rect 7350 61498 7356 61500
rect 7412 61498 7436 61500
rect 7492 61498 7516 61500
rect 7572 61498 7596 61500
rect 7652 61498 7658 61500
rect 7412 61446 7414 61498
rect 7594 61446 7596 61498
rect 7350 61444 7356 61446
rect 7412 61444 7436 61446
rect 7492 61444 7516 61446
rect 7572 61444 7596 61446
rect 7652 61444 7658 61446
rect 7350 61435 7658 61444
rect 7760 61282 7788 65350
rect 7852 65142 7880 65470
rect 7840 65136 7892 65142
rect 7840 65078 7892 65084
rect 7852 63578 7880 65078
rect 7944 64326 7972 65486
rect 8392 65408 8444 65414
rect 8392 65350 8444 65356
rect 8010 65308 8318 65317
rect 8010 65306 8016 65308
rect 8072 65306 8096 65308
rect 8152 65306 8176 65308
rect 8232 65306 8256 65308
rect 8312 65306 8318 65308
rect 8072 65254 8074 65306
rect 8254 65254 8256 65306
rect 8010 65252 8016 65254
rect 8072 65252 8096 65254
rect 8152 65252 8176 65254
rect 8232 65252 8256 65254
rect 8312 65252 8318 65254
rect 8010 65243 8318 65252
rect 8404 65113 8432 65350
rect 8390 65104 8446 65113
rect 8390 65039 8446 65048
rect 8208 64864 8260 64870
rect 8208 64806 8260 64812
rect 8220 64530 8248 64806
rect 8208 64524 8260 64530
rect 8208 64466 8260 64472
rect 7932 64320 7984 64326
rect 7932 64262 7984 64268
rect 7840 63572 7892 63578
rect 7840 63514 7892 63520
rect 7840 63436 7892 63442
rect 7840 63378 7892 63384
rect 7852 63050 7880 63378
rect 7944 63306 7972 64262
rect 8010 64220 8318 64229
rect 8010 64218 8016 64220
rect 8072 64218 8096 64220
rect 8152 64218 8176 64220
rect 8232 64218 8256 64220
rect 8312 64218 8318 64220
rect 8072 64166 8074 64218
rect 8254 64166 8256 64218
rect 8010 64164 8016 64166
rect 8072 64164 8096 64166
rect 8152 64164 8176 64166
rect 8232 64164 8256 64166
rect 8312 64164 8318 64166
rect 8010 64155 8318 64164
rect 8208 63776 8260 63782
rect 8208 63718 8260 63724
rect 8482 63744 8538 63753
rect 8220 63374 8248 63718
rect 8482 63679 8538 63688
rect 8496 63578 8524 63679
rect 8484 63572 8536 63578
rect 8484 63514 8536 63520
rect 8208 63368 8260 63374
rect 8208 63310 8260 63316
rect 7932 63300 7984 63306
rect 7932 63242 7984 63248
rect 8010 63132 8318 63141
rect 8010 63130 8016 63132
rect 8072 63130 8096 63132
rect 8152 63130 8176 63132
rect 8232 63130 8256 63132
rect 8312 63130 8318 63132
rect 8072 63078 8074 63130
rect 8254 63078 8256 63130
rect 8010 63076 8016 63078
rect 8072 63076 8096 63078
rect 8152 63076 8176 63078
rect 8232 63076 8256 63078
rect 8312 63076 8318 63078
rect 8010 63067 8318 63076
rect 7852 63022 7972 63050
rect 7300 61254 7788 61282
rect 7300 60734 7328 61254
rect 7748 61192 7800 61198
rect 7748 61134 7800 61140
rect 7380 61056 7432 61062
rect 7380 60998 7432 61004
rect 7392 60858 7420 60998
rect 7380 60852 7432 60858
rect 7380 60794 7432 60800
rect 7300 60706 7420 60734
rect 7392 60654 7420 60706
rect 7380 60648 7432 60654
rect 7380 60590 7432 60596
rect 7760 60518 7788 61134
rect 7944 61130 7972 63022
rect 8024 62892 8076 62898
rect 8024 62834 8076 62840
rect 8036 62150 8064 62834
rect 8392 62688 8444 62694
rect 8392 62630 8444 62636
rect 8404 62393 8432 62630
rect 8390 62384 8446 62393
rect 8390 62319 8446 62328
rect 8024 62144 8076 62150
rect 8024 62086 8076 62092
rect 8010 62044 8318 62053
rect 8010 62042 8016 62044
rect 8072 62042 8096 62044
rect 8152 62042 8176 62044
rect 8232 62042 8256 62044
rect 8312 62042 8318 62044
rect 8072 61990 8074 62042
rect 8254 61990 8256 62042
rect 8010 61988 8016 61990
rect 8072 61988 8096 61990
rect 8152 61988 8176 61990
rect 8232 61988 8256 61990
rect 8312 61988 8318 61990
rect 8010 61979 8318 61988
rect 7932 61124 7984 61130
rect 7932 61066 7984 61072
rect 7838 60616 7894 60625
rect 7838 60551 7894 60560
rect 7748 60512 7800 60518
rect 7748 60454 7800 60460
rect 7350 60412 7658 60421
rect 7350 60410 7356 60412
rect 7412 60410 7436 60412
rect 7492 60410 7516 60412
rect 7572 60410 7596 60412
rect 7652 60410 7658 60412
rect 7412 60358 7414 60410
rect 7594 60358 7596 60410
rect 7350 60356 7356 60358
rect 7412 60356 7436 60358
rect 7492 60356 7516 60358
rect 7572 60356 7596 60358
rect 7652 60356 7658 60358
rect 7350 60347 7658 60356
rect 7748 60104 7800 60110
rect 7748 60046 7800 60052
rect 7760 59430 7788 60046
rect 7748 59424 7800 59430
rect 7748 59366 7800 59372
rect 7350 59324 7658 59333
rect 7350 59322 7356 59324
rect 7412 59322 7436 59324
rect 7492 59322 7516 59324
rect 7572 59322 7596 59324
rect 7652 59322 7658 59324
rect 7412 59270 7414 59322
rect 7594 59270 7596 59322
rect 7350 59268 7356 59270
rect 7412 59268 7436 59270
rect 7492 59268 7516 59270
rect 7572 59268 7596 59270
rect 7652 59268 7658 59270
rect 7350 59259 7658 59268
rect 7748 58948 7800 58954
rect 7748 58890 7800 58896
rect 7760 58342 7788 58890
rect 7748 58336 7800 58342
rect 7748 58278 7800 58284
rect 7350 58236 7658 58245
rect 7350 58234 7356 58236
rect 7412 58234 7436 58236
rect 7492 58234 7516 58236
rect 7572 58234 7596 58236
rect 7652 58234 7658 58236
rect 7412 58182 7414 58234
rect 7594 58182 7596 58234
rect 7350 58180 7356 58182
rect 7412 58180 7436 58182
rect 7492 58180 7516 58182
rect 7572 58180 7596 58182
rect 7652 58180 7658 58182
rect 7350 58171 7658 58180
rect 7748 57996 7800 58002
rect 7748 57938 7800 57944
rect 7656 57792 7708 57798
rect 7656 57734 7708 57740
rect 7668 57390 7696 57734
rect 7656 57384 7708 57390
rect 7656 57326 7708 57332
rect 7350 57148 7658 57157
rect 7350 57146 7356 57148
rect 7412 57146 7436 57148
rect 7492 57146 7516 57148
rect 7572 57146 7596 57148
rect 7652 57146 7658 57148
rect 7412 57094 7414 57146
rect 7594 57094 7596 57146
rect 7350 57092 7356 57094
rect 7412 57092 7436 57094
rect 7492 57092 7516 57094
rect 7572 57092 7596 57094
rect 7652 57092 7658 57094
rect 7350 57083 7658 57092
rect 7656 56704 7708 56710
rect 7656 56646 7708 56652
rect 7668 56166 7696 56646
rect 7760 56302 7788 57938
rect 7748 56296 7800 56302
rect 7748 56238 7800 56244
rect 7656 56160 7708 56166
rect 7656 56102 7708 56108
rect 7350 56060 7658 56069
rect 7350 56058 7356 56060
rect 7412 56058 7436 56060
rect 7492 56058 7516 56060
rect 7572 56058 7596 56060
rect 7652 56058 7658 56060
rect 7412 56006 7414 56058
rect 7594 56006 7596 56058
rect 7350 56004 7356 56006
rect 7412 56004 7436 56006
rect 7492 56004 7516 56006
rect 7572 56004 7596 56006
rect 7652 56004 7658 56006
rect 7350 55995 7658 56004
rect 7350 54972 7658 54981
rect 7350 54970 7356 54972
rect 7412 54970 7436 54972
rect 7492 54970 7516 54972
rect 7572 54970 7596 54972
rect 7652 54970 7658 54972
rect 7412 54918 7414 54970
rect 7594 54918 7596 54970
rect 7350 54916 7356 54918
rect 7412 54916 7436 54918
rect 7492 54916 7516 54918
rect 7572 54916 7596 54918
rect 7652 54916 7658 54918
rect 7350 54907 7658 54916
rect 7656 54800 7708 54806
rect 7656 54742 7708 54748
rect 7668 54262 7696 54742
rect 7656 54256 7708 54262
rect 7656 54198 7708 54204
rect 7668 54126 7696 54198
rect 7656 54120 7708 54126
rect 7656 54062 7708 54068
rect 7350 53884 7658 53893
rect 7350 53882 7356 53884
rect 7412 53882 7436 53884
rect 7492 53882 7516 53884
rect 7572 53882 7596 53884
rect 7652 53882 7658 53884
rect 7412 53830 7414 53882
rect 7594 53830 7596 53882
rect 7350 53828 7356 53830
rect 7412 53828 7436 53830
rect 7492 53828 7516 53830
rect 7572 53828 7596 53830
rect 7652 53828 7658 53830
rect 7350 53819 7658 53828
rect 7350 52796 7658 52805
rect 7350 52794 7356 52796
rect 7412 52794 7436 52796
rect 7492 52794 7516 52796
rect 7572 52794 7596 52796
rect 7652 52794 7658 52796
rect 7412 52742 7414 52794
rect 7594 52742 7596 52794
rect 7350 52740 7356 52742
rect 7412 52740 7436 52742
rect 7492 52740 7516 52742
rect 7572 52740 7596 52742
rect 7652 52740 7658 52742
rect 7350 52731 7658 52740
rect 7350 51708 7658 51717
rect 7350 51706 7356 51708
rect 7412 51706 7436 51708
rect 7492 51706 7516 51708
rect 7572 51706 7596 51708
rect 7652 51706 7658 51708
rect 7412 51654 7414 51706
rect 7594 51654 7596 51706
rect 7350 51652 7356 51654
rect 7412 51652 7436 51654
rect 7492 51652 7516 51654
rect 7572 51652 7596 51654
rect 7652 51652 7658 51654
rect 7350 51643 7658 51652
rect 7380 51604 7432 51610
rect 7380 51546 7432 51552
rect 7392 50726 7420 51546
rect 7852 50844 7880 60551
rect 7944 56234 7972 61066
rect 8392 61056 8444 61062
rect 8390 61024 8392 61033
rect 8444 61024 8446 61033
rect 8010 60956 8318 60965
rect 8390 60959 8446 60968
rect 8010 60954 8016 60956
rect 8072 60954 8096 60956
rect 8152 60954 8176 60956
rect 8232 60954 8256 60956
rect 8312 60954 8318 60956
rect 8072 60902 8074 60954
rect 8254 60902 8256 60954
rect 8010 60900 8016 60902
rect 8072 60900 8096 60902
rect 8152 60900 8176 60902
rect 8232 60900 8256 60902
rect 8312 60900 8318 60902
rect 8010 60891 8318 60900
rect 8024 60852 8076 60858
rect 8024 60794 8076 60800
rect 8036 60178 8064 60794
rect 8024 60172 8076 60178
rect 8024 60114 8076 60120
rect 8392 59968 8444 59974
rect 8392 59910 8444 59916
rect 8010 59868 8318 59877
rect 8010 59866 8016 59868
rect 8072 59866 8096 59868
rect 8152 59866 8176 59868
rect 8232 59866 8256 59868
rect 8312 59866 8318 59868
rect 8072 59814 8074 59866
rect 8254 59814 8256 59866
rect 8010 59812 8016 59814
rect 8072 59812 8096 59814
rect 8152 59812 8176 59814
rect 8232 59812 8256 59814
rect 8312 59812 8318 59814
rect 8010 59803 8318 59812
rect 8404 59673 8432 59910
rect 8390 59664 8446 59673
rect 8390 59599 8446 59608
rect 8484 58880 8536 58886
rect 8484 58822 8536 58828
rect 8010 58780 8318 58789
rect 8010 58778 8016 58780
rect 8072 58778 8096 58780
rect 8152 58778 8176 58780
rect 8232 58778 8256 58780
rect 8312 58778 8318 58780
rect 8072 58726 8074 58778
rect 8254 58726 8256 58778
rect 8010 58724 8016 58726
rect 8072 58724 8096 58726
rect 8152 58724 8176 58726
rect 8232 58724 8256 58726
rect 8312 58724 8318 58726
rect 8010 58715 8318 58724
rect 8496 58313 8524 58822
rect 8482 58304 8538 58313
rect 8482 58239 8538 58248
rect 8010 57692 8318 57701
rect 8010 57690 8016 57692
rect 8072 57690 8096 57692
rect 8152 57690 8176 57692
rect 8232 57690 8256 57692
rect 8312 57690 8318 57692
rect 8072 57638 8074 57690
rect 8254 57638 8256 57690
rect 8010 57636 8016 57638
rect 8072 57636 8096 57638
rect 8152 57636 8176 57638
rect 8232 57636 8256 57638
rect 8312 57636 8318 57638
rect 8010 57627 8318 57636
rect 8024 57384 8076 57390
rect 8024 57326 8076 57332
rect 8036 56846 8064 57326
rect 8576 57248 8628 57254
rect 8576 57190 8628 57196
rect 8588 56953 8616 57190
rect 8574 56944 8630 56953
rect 8574 56879 8630 56888
rect 8024 56840 8076 56846
rect 8024 56782 8076 56788
rect 8010 56604 8318 56613
rect 8010 56602 8016 56604
rect 8072 56602 8096 56604
rect 8152 56602 8176 56604
rect 8232 56602 8256 56604
rect 8312 56602 8318 56604
rect 8072 56550 8074 56602
rect 8254 56550 8256 56602
rect 8010 56548 8016 56550
rect 8072 56548 8096 56550
rect 8152 56548 8176 56550
rect 8232 56548 8256 56550
rect 8312 56548 8318 56550
rect 8010 56539 8318 56548
rect 7932 56228 7984 56234
rect 7932 56170 7984 56176
rect 8024 56160 8076 56166
rect 8024 56102 8076 56108
rect 8036 55758 8064 56102
rect 8024 55752 8076 55758
rect 7944 55700 8024 55706
rect 7944 55694 8076 55700
rect 7944 55678 8064 55694
rect 7944 54806 7972 55678
rect 8484 55616 8536 55622
rect 8484 55558 8536 55564
rect 8010 55516 8318 55525
rect 8010 55514 8016 55516
rect 8072 55514 8096 55516
rect 8152 55514 8176 55516
rect 8232 55514 8256 55516
rect 8312 55514 8318 55516
rect 8072 55462 8074 55514
rect 8254 55462 8256 55514
rect 8010 55460 8016 55462
rect 8072 55460 8096 55462
rect 8152 55460 8176 55462
rect 8232 55460 8256 55462
rect 8312 55460 8318 55462
rect 8010 55451 8318 55460
rect 8206 55312 8262 55321
rect 8496 55282 8524 55558
rect 8206 55247 8262 55256
rect 8484 55276 8536 55282
rect 8220 54874 8248 55247
rect 8484 55218 8536 55224
rect 8208 54868 8260 54874
rect 8208 54810 8260 54816
rect 7932 54800 7984 54806
rect 7932 54742 7984 54748
rect 8496 54670 8524 55218
rect 7932 54664 7984 54670
rect 7932 54606 7984 54612
rect 8484 54664 8536 54670
rect 8484 54606 8536 54612
rect 7944 54210 7972 54606
rect 8392 54528 8444 54534
rect 8392 54470 8444 54476
rect 8010 54428 8318 54437
rect 8010 54426 8016 54428
rect 8072 54426 8096 54428
rect 8152 54426 8176 54428
rect 8232 54426 8256 54428
rect 8312 54426 8318 54428
rect 8072 54374 8074 54426
rect 8254 54374 8256 54426
rect 8010 54372 8016 54374
rect 8072 54372 8096 54374
rect 8152 54372 8176 54374
rect 8232 54372 8256 54374
rect 8312 54372 8318 54374
rect 8010 54363 8318 54372
rect 8404 54233 8432 54470
rect 8390 54224 8446 54233
rect 7944 54182 8064 54210
rect 8036 53990 8064 54182
rect 8390 54159 8446 54168
rect 8116 54052 8168 54058
rect 8116 53994 8168 54000
rect 8024 53984 8076 53990
rect 8024 53926 8076 53932
rect 8128 53802 8156 53994
rect 7944 53774 8156 53802
rect 7944 53242 7972 53774
rect 8010 53340 8318 53349
rect 8010 53338 8016 53340
rect 8072 53338 8096 53340
rect 8152 53338 8176 53340
rect 8232 53338 8256 53340
rect 8312 53338 8318 53340
rect 8072 53286 8074 53338
rect 8254 53286 8256 53338
rect 8010 53284 8016 53286
rect 8072 53284 8096 53286
rect 8152 53284 8176 53286
rect 8232 53284 8256 53286
rect 8312 53284 8318 53286
rect 8010 53275 8318 53284
rect 7932 53236 7984 53242
rect 7932 53178 7984 53184
rect 7944 52154 7972 53178
rect 8208 52896 8260 52902
rect 8208 52838 8260 52844
rect 8390 52864 8446 52873
rect 8220 52494 8248 52838
rect 8390 52799 8446 52808
rect 8404 52698 8432 52799
rect 8392 52692 8444 52698
rect 8392 52634 8444 52640
rect 8208 52488 8260 52494
rect 8208 52430 8260 52436
rect 8010 52252 8318 52261
rect 8010 52250 8016 52252
rect 8072 52250 8096 52252
rect 8152 52250 8176 52252
rect 8232 52250 8256 52252
rect 8312 52250 8318 52252
rect 8072 52198 8074 52250
rect 8254 52198 8256 52250
rect 8010 52196 8016 52198
rect 8072 52196 8096 52198
rect 8152 52196 8176 52198
rect 8232 52196 8256 52198
rect 8312 52196 8318 52198
rect 8010 52187 8318 52196
rect 7932 52148 7984 52154
rect 7932 52090 7984 52096
rect 8116 52148 8168 52154
rect 8116 52090 8168 52096
rect 7932 52012 7984 52018
rect 7932 51954 7984 51960
rect 7944 51270 7972 51954
rect 8128 51406 8156 52090
rect 8392 51808 8444 51814
rect 8392 51750 8444 51756
rect 8404 51513 8432 51750
rect 8390 51504 8446 51513
rect 8390 51439 8446 51448
rect 8116 51400 8168 51406
rect 8116 51342 8168 51348
rect 7932 51264 7984 51270
rect 7932 51206 7984 51212
rect 7944 51066 7972 51206
rect 8010 51164 8318 51173
rect 8010 51162 8016 51164
rect 8072 51162 8096 51164
rect 8152 51162 8176 51164
rect 8232 51162 8256 51164
rect 8312 51162 8318 51164
rect 8072 51110 8074 51162
rect 8254 51110 8256 51162
rect 8010 51108 8016 51110
rect 8072 51108 8096 51110
rect 8152 51108 8176 51110
rect 8232 51108 8256 51110
rect 8312 51108 8318 51110
rect 8010 51099 8318 51108
rect 7932 51060 7984 51066
rect 7932 51002 7984 51008
rect 7760 50816 7880 50844
rect 7380 50720 7432 50726
rect 7380 50662 7432 50668
rect 7350 50620 7658 50629
rect 7350 50618 7356 50620
rect 7412 50618 7436 50620
rect 7492 50618 7516 50620
rect 7572 50618 7596 50620
rect 7652 50618 7658 50620
rect 7412 50566 7414 50618
rect 7594 50566 7596 50618
rect 7350 50564 7356 50566
rect 7412 50564 7436 50566
rect 7492 50564 7516 50566
rect 7572 50564 7596 50566
rect 7652 50564 7658 50566
rect 7350 50555 7658 50564
rect 7350 49532 7658 49541
rect 7350 49530 7356 49532
rect 7412 49530 7436 49532
rect 7492 49530 7516 49532
rect 7572 49530 7596 49532
rect 7652 49530 7658 49532
rect 7412 49478 7414 49530
rect 7594 49478 7596 49530
rect 7350 49476 7356 49478
rect 7412 49476 7436 49478
rect 7492 49476 7516 49478
rect 7572 49476 7596 49478
rect 7652 49476 7658 49478
rect 7350 49467 7658 49476
rect 7472 49428 7524 49434
rect 7472 49370 7524 49376
rect 7288 49088 7340 49094
rect 7288 49030 7340 49036
rect 7300 48890 7328 49030
rect 7288 48884 7340 48890
rect 7288 48826 7340 48832
rect 7484 48822 7512 49370
rect 7760 49314 7788 50816
rect 7840 50720 7892 50726
rect 7840 50662 7892 50668
rect 7668 49286 7788 49314
rect 7472 48816 7524 48822
rect 7472 48758 7524 48764
rect 7668 48686 7696 49286
rect 7748 49224 7800 49230
rect 7748 49166 7800 49172
rect 7656 48680 7708 48686
rect 7656 48622 7708 48628
rect 7350 48444 7658 48453
rect 7350 48442 7356 48444
rect 7412 48442 7436 48444
rect 7492 48442 7516 48444
rect 7572 48442 7596 48444
rect 7652 48442 7658 48444
rect 7412 48390 7414 48442
rect 7594 48390 7596 48442
rect 7350 48388 7356 48390
rect 7412 48388 7436 48390
rect 7492 48388 7516 48390
rect 7572 48388 7596 48390
rect 7652 48388 7658 48390
rect 7350 48379 7658 48388
rect 7760 48346 7788 49166
rect 7748 48340 7800 48346
rect 7748 48282 7800 48288
rect 7852 48226 7880 50662
rect 7932 50176 7984 50182
rect 7932 50118 7984 50124
rect 8390 50144 8446 50153
rect 7944 49434 7972 50118
rect 8010 50076 8318 50085
rect 8390 50079 8446 50088
rect 8010 50074 8016 50076
rect 8072 50074 8096 50076
rect 8152 50074 8176 50076
rect 8232 50074 8256 50076
rect 8312 50074 8318 50076
rect 8072 50022 8074 50074
rect 8254 50022 8256 50074
rect 8010 50020 8016 50022
rect 8072 50020 8096 50022
rect 8152 50020 8176 50022
rect 8232 50020 8256 50022
rect 8312 50020 8318 50022
rect 8010 50011 8318 50020
rect 8404 49978 8432 50079
rect 8392 49972 8444 49978
rect 8392 49914 8444 49920
rect 7932 49428 7984 49434
rect 7932 49370 7984 49376
rect 7932 49224 7984 49230
rect 7932 49166 7984 49172
rect 7944 48770 7972 49166
rect 8392 49088 8444 49094
rect 8392 49030 8444 49036
rect 8010 48988 8318 48997
rect 8010 48986 8016 48988
rect 8072 48986 8096 48988
rect 8152 48986 8176 48988
rect 8232 48986 8256 48988
rect 8312 48986 8318 48988
rect 8072 48934 8074 48986
rect 8254 48934 8256 48986
rect 8010 48932 8016 48934
rect 8072 48932 8096 48934
rect 8152 48932 8176 48934
rect 8232 48932 8256 48934
rect 8312 48932 8318 48934
rect 8010 48923 8318 48932
rect 8404 48793 8432 49030
rect 8390 48784 8446 48793
rect 7944 48742 8064 48770
rect 8036 48550 8064 48742
rect 8390 48719 8446 48728
rect 8024 48544 8076 48550
rect 8024 48486 8076 48492
rect 7760 48198 7880 48226
rect 7350 47356 7658 47365
rect 7350 47354 7356 47356
rect 7412 47354 7436 47356
rect 7492 47354 7516 47356
rect 7572 47354 7596 47356
rect 7652 47354 7658 47356
rect 7412 47302 7414 47354
rect 7594 47302 7596 47354
rect 7350 47300 7356 47302
rect 7412 47300 7436 47302
rect 7492 47300 7516 47302
rect 7572 47300 7596 47302
rect 7652 47300 7658 47302
rect 7350 47291 7658 47300
rect 7380 47116 7432 47122
rect 7380 47058 7432 47064
rect 7392 46510 7420 47058
rect 7380 46504 7432 46510
rect 7380 46446 7432 46452
rect 7350 46268 7658 46277
rect 7350 46266 7356 46268
rect 7412 46266 7436 46268
rect 7492 46266 7516 46268
rect 7572 46266 7596 46268
rect 7652 46266 7658 46268
rect 7412 46214 7414 46266
rect 7594 46214 7596 46266
rect 7350 46212 7356 46214
rect 7412 46212 7436 46214
rect 7492 46212 7516 46214
rect 7572 46212 7596 46214
rect 7652 46212 7658 46214
rect 7350 46203 7658 46212
rect 7024 45614 7236 45642
rect 6920 45484 6972 45490
rect 6920 45426 6972 45432
rect 6920 45280 6972 45286
rect 6920 45222 6972 45228
rect 6932 44538 6960 45222
rect 6920 44532 6972 44538
rect 6920 44474 6972 44480
rect 6920 43444 6972 43450
rect 6920 43386 6972 43392
rect 6932 43194 6960 43386
rect 6840 43166 6960 43194
rect 6840 42786 6868 43166
rect 6920 43104 6972 43110
rect 6920 43046 6972 43052
rect 6932 42906 6960 43046
rect 6920 42900 6972 42906
rect 6920 42842 6972 42848
rect 6840 42758 6960 42786
rect 6828 42628 6880 42634
rect 6828 42570 6880 42576
rect 6736 41608 6788 41614
rect 6736 41550 6788 41556
rect 6840 41414 6868 42570
rect 6932 42158 6960 42758
rect 6920 42152 6972 42158
rect 6920 42094 6972 42100
rect 6932 41614 6960 42094
rect 6920 41608 6972 41614
rect 6920 41550 6972 41556
rect 6840 41386 6960 41414
rect 6932 41206 6960 41386
rect 6920 41200 6972 41206
rect 6920 41142 6972 41148
rect 6460 41132 6512 41138
rect 6460 41074 6512 41080
rect 6472 40186 6500 41074
rect 6920 40928 6972 40934
rect 6920 40870 6972 40876
rect 6736 40520 6788 40526
rect 6736 40462 6788 40468
rect 6092 40180 6144 40186
rect 6092 40122 6144 40128
rect 6368 40180 6420 40186
rect 6368 40122 6420 40128
rect 6460 40180 6512 40186
rect 6460 40122 6512 40128
rect 5908 39976 5960 39982
rect 5908 39918 5960 39924
rect 6276 39976 6328 39982
rect 6276 39918 6328 39924
rect 2350 39740 2658 39749
rect 2350 39738 2356 39740
rect 2412 39738 2436 39740
rect 2492 39738 2516 39740
rect 2572 39738 2596 39740
rect 2652 39738 2658 39740
rect 2412 39686 2414 39738
rect 2594 39686 2596 39738
rect 2350 39684 2356 39686
rect 2412 39684 2436 39686
rect 2492 39684 2516 39686
rect 2572 39684 2596 39686
rect 2652 39684 2658 39686
rect 2350 39675 2658 39684
rect 4436 39432 4488 39438
rect 4436 39374 4488 39380
rect 3010 39196 3318 39205
rect 3010 39194 3016 39196
rect 3072 39194 3096 39196
rect 3152 39194 3176 39196
rect 3232 39194 3256 39196
rect 3312 39194 3318 39196
rect 3072 39142 3074 39194
rect 3254 39142 3256 39194
rect 3010 39140 3016 39142
rect 3072 39140 3096 39142
rect 3152 39140 3176 39142
rect 3232 39140 3256 39142
rect 3312 39140 3318 39142
rect 3010 39131 3318 39140
rect 2350 38652 2658 38661
rect 2350 38650 2356 38652
rect 2412 38650 2436 38652
rect 2492 38650 2516 38652
rect 2572 38650 2596 38652
rect 2652 38650 2658 38652
rect 2412 38598 2414 38650
rect 2594 38598 2596 38650
rect 2350 38596 2356 38598
rect 2412 38596 2436 38598
rect 2492 38596 2516 38598
rect 2572 38596 2596 38598
rect 2652 38596 2658 38598
rect 2350 38587 2658 38596
rect 4448 38350 4476 39374
rect 4988 39364 5040 39370
rect 4988 39306 5040 39312
rect 5000 39098 5028 39306
rect 5908 39296 5960 39302
rect 5908 39238 5960 39244
rect 4988 39092 5040 39098
rect 4988 39034 5040 39040
rect 5920 38962 5948 39238
rect 6288 39030 6316 39918
rect 6552 39840 6604 39846
rect 6552 39782 6604 39788
rect 6564 39370 6592 39782
rect 6748 39438 6776 40462
rect 6932 40458 6960 40870
rect 7024 40594 7052 45614
rect 7104 45484 7156 45490
rect 7104 45426 7156 45432
rect 7116 43450 7144 45426
rect 7350 45180 7658 45189
rect 7350 45178 7356 45180
rect 7412 45178 7436 45180
rect 7492 45178 7516 45180
rect 7572 45178 7596 45180
rect 7652 45178 7658 45180
rect 7412 45126 7414 45178
rect 7594 45126 7596 45178
rect 7350 45124 7356 45126
rect 7412 45124 7436 45126
rect 7492 45124 7516 45126
rect 7572 45124 7596 45126
rect 7652 45124 7658 45126
rect 7350 45115 7658 45124
rect 7196 44736 7248 44742
rect 7196 44678 7248 44684
rect 7208 44538 7236 44678
rect 7196 44532 7248 44538
rect 7196 44474 7248 44480
rect 7350 44092 7658 44101
rect 7350 44090 7356 44092
rect 7412 44090 7436 44092
rect 7492 44090 7516 44092
rect 7572 44090 7596 44092
rect 7652 44090 7658 44092
rect 7412 44038 7414 44090
rect 7594 44038 7596 44090
rect 7350 44036 7356 44038
rect 7412 44036 7436 44038
rect 7492 44036 7516 44038
rect 7572 44036 7596 44038
rect 7652 44036 7658 44038
rect 7350 44027 7658 44036
rect 7104 43444 7156 43450
rect 7104 43386 7156 43392
rect 7104 43308 7156 43314
rect 7104 43250 7156 43256
rect 7196 43308 7248 43314
rect 7196 43250 7248 43256
rect 7116 42566 7144 43250
rect 7104 42560 7156 42566
rect 7104 42502 7156 42508
rect 7116 42362 7144 42502
rect 7208 42362 7236 43250
rect 7350 43004 7658 43013
rect 7350 43002 7356 43004
rect 7412 43002 7436 43004
rect 7492 43002 7516 43004
rect 7572 43002 7596 43004
rect 7652 43002 7658 43004
rect 7412 42950 7414 43002
rect 7594 42950 7596 43002
rect 7350 42948 7356 42950
rect 7412 42948 7436 42950
rect 7492 42948 7516 42950
rect 7572 42948 7596 42950
rect 7652 42948 7658 42950
rect 7350 42939 7658 42948
rect 7104 42356 7156 42362
rect 7104 42298 7156 42304
rect 7196 42356 7248 42362
rect 7196 42298 7248 42304
rect 7760 42242 7788 48198
rect 8036 48142 8064 48486
rect 8024 48136 8076 48142
rect 8024 48078 8076 48084
rect 8010 47900 8318 47909
rect 8010 47898 8016 47900
rect 8072 47898 8096 47900
rect 8152 47898 8176 47900
rect 8232 47898 8256 47900
rect 8312 47898 8318 47900
rect 8072 47846 8074 47898
rect 8254 47846 8256 47898
rect 8010 47844 8016 47846
rect 8072 47844 8096 47846
rect 8152 47844 8176 47846
rect 8232 47844 8256 47846
rect 8312 47844 8318 47846
rect 8010 47835 8318 47844
rect 8390 47424 8446 47433
rect 8390 47359 8446 47368
rect 8404 47258 8432 47359
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 8010 46812 8318 46821
rect 8010 46810 8016 46812
rect 8072 46810 8096 46812
rect 8152 46810 8176 46812
rect 8232 46810 8256 46812
rect 8312 46810 8318 46812
rect 8072 46758 8074 46810
rect 8254 46758 8256 46810
rect 8010 46756 8016 46758
rect 8072 46756 8096 46758
rect 8152 46756 8176 46758
rect 8232 46756 8256 46758
rect 8312 46756 8318 46758
rect 8010 46747 8318 46756
rect 8024 46640 8076 46646
rect 8024 46582 8076 46588
rect 7840 46504 7892 46510
rect 7840 46446 7892 46452
rect 7852 45422 7880 46446
rect 8036 45966 8064 46582
rect 8392 46368 8444 46374
rect 8392 46310 8444 46316
rect 8404 46073 8432 46310
rect 8390 46064 8446 46073
rect 8390 45999 8446 46008
rect 8024 45960 8076 45966
rect 7944 45908 8024 45914
rect 7944 45902 8076 45908
rect 7944 45886 8064 45902
rect 7840 45416 7892 45422
rect 7840 45358 7892 45364
rect 7944 44962 7972 45886
rect 8010 45724 8318 45733
rect 8010 45722 8016 45724
rect 8072 45722 8096 45724
rect 8152 45722 8176 45724
rect 8232 45722 8256 45724
rect 8312 45722 8318 45724
rect 8072 45670 8074 45722
rect 8254 45670 8256 45722
rect 8010 45668 8016 45670
rect 8072 45668 8096 45670
rect 8152 45668 8176 45670
rect 8232 45668 8256 45670
rect 8312 45668 8318 45670
rect 8010 45659 8318 45668
rect 7944 44934 8064 44962
rect 8036 44878 8064 44934
rect 8024 44872 8076 44878
rect 8024 44814 8076 44820
rect 8390 44704 8446 44713
rect 8010 44636 8318 44645
rect 8390 44639 8446 44648
rect 8010 44634 8016 44636
rect 8072 44634 8096 44636
rect 8152 44634 8176 44636
rect 8232 44634 8256 44636
rect 8312 44634 8318 44636
rect 8072 44582 8074 44634
rect 8254 44582 8256 44634
rect 8010 44580 8016 44582
rect 8072 44580 8096 44582
rect 8152 44580 8176 44582
rect 8232 44580 8256 44582
rect 8312 44580 8318 44582
rect 8010 44571 8318 44580
rect 8404 44538 8432 44639
rect 8392 44532 8444 44538
rect 8392 44474 8444 44480
rect 7932 43648 7984 43654
rect 7932 43590 7984 43596
rect 8852 43648 8904 43654
rect 8852 43590 8904 43596
rect 7840 42560 7892 42566
rect 7840 42502 7892 42508
rect 7852 42294 7880 42502
rect 7944 42294 7972 43590
rect 8010 43548 8318 43557
rect 8010 43546 8016 43548
rect 8072 43546 8096 43548
rect 8152 43546 8176 43548
rect 8232 43546 8256 43548
rect 8312 43546 8318 43548
rect 8072 43494 8074 43546
rect 8254 43494 8256 43546
rect 8010 43492 8016 43494
rect 8072 43492 8096 43494
rect 8152 43492 8176 43494
rect 8232 43492 8256 43494
rect 8312 43492 8318 43494
rect 8010 43483 8318 43492
rect 8864 43353 8892 43590
rect 8850 43344 8906 43353
rect 8850 43279 8906 43288
rect 8010 42460 8318 42469
rect 8010 42458 8016 42460
rect 8072 42458 8096 42460
rect 8152 42458 8176 42460
rect 8232 42458 8256 42460
rect 8312 42458 8318 42460
rect 8072 42406 8074 42458
rect 8254 42406 8256 42458
rect 8010 42404 8016 42406
rect 8072 42404 8096 42406
rect 8152 42404 8176 42406
rect 8232 42404 8256 42406
rect 8312 42404 8318 42406
rect 8010 42395 8318 42404
rect 7208 42214 7788 42242
rect 7840 42288 7892 42294
rect 7840 42230 7892 42236
rect 7932 42288 7984 42294
rect 7932 42230 7984 42236
rect 7104 41200 7156 41206
rect 7104 41142 7156 41148
rect 7012 40588 7064 40594
rect 7012 40530 7064 40536
rect 7116 40458 7144 41142
rect 6920 40452 6972 40458
rect 6920 40394 6972 40400
rect 7104 40452 7156 40458
rect 7104 40394 7156 40400
rect 6828 40384 6880 40390
rect 7208 40338 7236 42214
rect 8392 42084 8444 42090
rect 8392 42026 8444 42032
rect 8404 41993 8432 42026
rect 8390 41984 8446 41993
rect 7350 41916 7658 41925
rect 8390 41919 8446 41928
rect 7350 41914 7356 41916
rect 7412 41914 7436 41916
rect 7492 41914 7516 41916
rect 7572 41914 7596 41916
rect 7652 41914 7658 41916
rect 7412 41862 7414 41914
rect 7594 41862 7596 41914
rect 7350 41860 7356 41862
rect 7412 41860 7436 41862
rect 7492 41860 7516 41862
rect 7572 41860 7596 41862
rect 7652 41860 7658 41862
rect 7350 41851 7658 41860
rect 7840 41540 7892 41546
rect 7840 41482 7892 41488
rect 7748 41472 7800 41478
rect 7748 41414 7800 41420
rect 7350 40828 7658 40837
rect 7350 40826 7356 40828
rect 7412 40826 7436 40828
rect 7492 40826 7516 40828
rect 7572 40826 7596 40828
rect 7652 40826 7658 40828
rect 7412 40774 7414 40826
rect 7594 40774 7596 40826
rect 7350 40772 7356 40774
rect 7412 40772 7436 40774
rect 7492 40772 7516 40774
rect 7572 40772 7596 40774
rect 7652 40772 7658 40774
rect 7350 40763 7658 40772
rect 6828 40326 6880 40332
rect 6736 39432 6788 39438
rect 6736 39374 6788 39380
rect 6552 39364 6604 39370
rect 6552 39306 6604 39312
rect 6276 39024 6328 39030
rect 6276 38966 6328 38972
rect 5908 38956 5960 38962
rect 5908 38898 5960 38904
rect 4436 38344 4488 38350
rect 4436 38286 4488 38292
rect 3010 38108 3318 38117
rect 3010 38106 3016 38108
rect 3072 38106 3096 38108
rect 3152 38106 3176 38108
rect 3232 38106 3256 38108
rect 3312 38106 3318 38108
rect 3072 38054 3074 38106
rect 3254 38054 3256 38106
rect 3010 38052 3016 38054
rect 3072 38052 3096 38054
rect 3152 38052 3176 38054
rect 3232 38052 3256 38054
rect 3312 38052 3318 38054
rect 3010 38043 3318 38052
rect 2350 37564 2658 37573
rect 2350 37562 2356 37564
rect 2412 37562 2436 37564
rect 2492 37562 2516 37564
rect 2572 37562 2596 37564
rect 2652 37562 2658 37564
rect 2412 37510 2414 37562
rect 2594 37510 2596 37562
rect 2350 37508 2356 37510
rect 2412 37508 2436 37510
rect 2492 37508 2516 37510
rect 2572 37508 2596 37510
rect 2652 37508 2658 37510
rect 2350 37499 2658 37508
rect 3010 37020 3318 37029
rect 3010 37018 3016 37020
rect 3072 37018 3096 37020
rect 3152 37018 3176 37020
rect 3232 37018 3256 37020
rect 3312 37018 3318 37020
rect 3072 36966 3074 37018
rect 3254 36966 3256 37018
rect 3010 36964 3016 36966
rect 3072 36964 3096 36966
rect 3152 36964 3176 36966
rect 3232 36964 3256 36966
rect 3312 36964 3318 36966
rect 3010 36955 3318 36964
rect 4448 36718 4476 38286
rect 4896 38276 4948 38282
rect 4896 38218 4948 38224
rect 4908 38010 4936 38218
rect 5816 38208 5868 38214
rect 5816 38150 5868 38156
rect 4896 38004 4948 38010
rect 4896 37946 4948 37952
rect 5828 37890 5856 38150
rect 5920 38010 5948 38898
rect 6092 38888 6144 38894
rect 6092 38830 6144 38836
rect 6000 38344 6052 38350
rect 6000 38286 6052 38292
rect 5908 38004 5960 38010
rect 5908 37946 5960 37952
rect 5828 37862 5948 37890
rect 5920 37806 5948 37862
rect 5908 37800 5960 37806
rect 5908 37742 5960 37748
rect 5920 37194 5948 37742
rect 5908 37188 5960 37194
rect 5908 37130 5960 37136
rect 5080 37120 5132 37126
rect 5080 37062 5132 37068
rect 5092 36922 5120 37062
rect 5080 36916 5132 36922
rect 5080 36858 5132 36864
rect 4436 36712 4488 36718
rect 4436 36654 4488 36660
rect 2350 36476 2658 36485
rect 2350 36474 2356 36476
rect 2412 36474 2436 36476
rect 2492 36474 2516 36476
rect 2572 36474 2596 36476
rect 2652 36474 2658 36476
rect 2412 36422 2414 36474
rect 2594 36422 2596 36474
rect 2350 36420 2356 36422
rect 2412 36420 2436 36422
rect 2492 36420 2516 36422
rect 2572 36420 2596 36422
rect 2652 36420 2658 36422
rect 2350 36411 2658 36420
rect 3010 35932 3318 35941
rect 3010 35930 3016 35932
rect 3072 35930 3096 35932
rect 3152 35930 3176 35932
rect 3232 35930 3256 35932
rect 3312 35930 3318 35932
rect 3072 35878 3074 35930
rect 3254 35878 3256 35930
rect 3010 35876 3016 35878
rect 3072 35876 3096 35878
rect 3152 35876 3176 35878
rect 3232 35876 3256 35878
rect 3312 35876 3318 35878
rect 3010 35867 3318 35876
rect 2350 35388 2658 35397
rect 2350 35386 2356 35388
rect 2412 35386 2436 35388
rect 2492 35386 2516 35388
rect 2572 35386 2596 35388
rect 2652 35386 2658 35388
rect 2412 35334 2414 35386
rect 2594 35334 2596 35386
rect 2350 35332 2356 35334
rect 2412 35332 2436 35334
rect 2492 35332 2516 35334
rect 2572 35332 2596 35334
rect 2652 35332 2658 35334
rect 2350 35323 2658 35332
rect 4448 35086 4476 36654
rect 6012 36650 6040 38286
rect 6104 37806 6132 38830
rect 6092 37800 6144 37806
rect 6092 37742 6144 37748
rect 6104 37330 6132 37742
rect 6092 37324 6144 37330
rect 6092 37266 6144 37272
rect 6000 36644 6052 36650
rect 6000 36586 6052 36592
rect 6104 35894 6132 37266
rect 6184 37120 6236 37126
rect 6184 37062 6236 37068
rect 6196 36922 6224 37062
rect 6184 36916 6236 36922
rect 6184 36858 6236 36864
rect 6196 36242 6224 36858
rect 6184 36236 6236 36242
rect 6184 36178 6236 36184
rect 6012 35866 6132 35894
rect 5908 35624 5960 35630
rect 5908 35566 5960 35572
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 5000 35154 5028 35430
rect 5920 35290 5948 35566
rect 5908 35284 5960 35290
rect 5908 35226 5960 35232
rect 4988 35148 5040 35154
rect 4988 35090 5040 35096
rect 4436 35080 4488 35086
rect 4436 35022 4488 35028
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 3010 34844 3318 34853
rect 3010 34842 3016 34844
rect 3072 34842 3096 34844
rect 3152 34842 3176 34844
rect 3232 34842 3256 34844
rect 3312 34842 3318 34844
rect 3072 34790 3074 34842
rect 3254 34790 3256 34842
rect 3010 34788 3016 34790
rect 3072 34788 3096 34790
rect 3152 34788 3176 34790
rect 3232 34788 3256 34790
rect 3312 34788 3318 34790
rect 3010 34779 3318 34788
rect 4816 34542 4844 34886
rect 5448 34604 5500 34610
rect 5448 34546 5500 34552
rect 4804 34536 4856 34542
rect 4804 34478 4856 34484
rect 2350 34300 2658 34309
rect 2350 34298 2356 34300
rect 2412 34298 2436 34300
rect 2492 34298 2516 34300
rect 2572 34298 2596 34300
rect 2652 34298 2658 34300
rect 2412 34246 2414 34298
rect 2594 34246 2596 34298
rect 2350 34244 2356 34246
rect 2412 34244 2436 34246
rect 2492 34244 2516 34246
rect 2572 34244 2596 34246
rect 2652 34244 2658 34246
rect 2350 34235 2658 34244
rect 4816 34134 4844 34478
rect 4804 34128 4856 34134
rect 4804 34070 4856 34076
rect 3010 33756 3318 33765
rect 3010 33754 3016 33756
rect 3072 33754 3096 33756
rect 3152 33754 3176 33756
rect 3232 33754 3256 33756
rect 3312 33754 3318 33756
rect 3072 33702 3074 33754
rect 3254 33702 3256 33754
rect 3010 33700 3016 33702
rect 3072 33700 3096 33702
rect 3152 33700 3176 33702
rect 3232 33700 3256 33702
rect 3312 33700 3318 33702
rect 3010 33691 3318 33700
rect 2350 33212 2658 33221
rect 2350 33210 2356 33212
rect 2412 33210 2436 33212
rect 2492 33210 2516 33212
rect 2572 33210 2596 33212
rect 2652 33210 2658 33212
rect 2412 33158 2414 33210
rect 2594 33158 2596 33210
rect 2350 33156 2356 33158
rect 2412 33156 2436 33158
rect 2492 33156 2516 33158
rect 2572 33156 2596 33158
rect 2652 33156 2658 33158
rect 2350 33147 2658 33156
rect 3010 32668 3318 32677
rect 3010 32666 3016 32668
rect 3072 32666 3096 32668
rect 3152 32666 3176 32668
rect 3232 32666 3256 32668
rect 3312 32666 3318 32668
rect 3072 32614 3074 32666
rect 3254 32614 3256 32666
rect 3010 32612 3016 32614
rect 3072 32612 3096 32614
rect 3152 32612 3176 32614
rect 3232 32612 3256 32614
rect 3312 32612 3318 32614
rect 3010 32603 3318 32612
rect 4712 32360 4764 32366
rect 4712 32302 4764 32308
rect 2350 32124 2658 32133
rect 2350 32122 2356 32124
rect 2412 32122 2436 32124
rect 2492 32122 2516 32124
rect 2572 32122 2596 32124
rect 2652 32122 2658 32124
rect 2412 32070 2414 32122
rect 2594 32070 2596 32122
rect 2350 32068 2356 32070
rect 2412 32068 2436 32070
rect 2492 32068 2516 32070
rect 2572 32068 2596 32070
rect 2652 32068 2658 32070
rect 2350 32059 2658 32068
rect 4724 32026 4752 32302
rect 4816 32230 4844 34070
rect 5460 33658 5488 34546
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 5644 34202 5672 34342
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 5816 33652 5868 33658
rect 5920 33640 5948 35226
rect 5868 33612 5948 33640
rect 5816 33594 5868 33600
rect 4804 32224 4856 32230
rect 4804 32166 4856 32172
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 3010 31580 3318 31589
rect 3010 31578 3016 31580
rect 3072 31578 3096 31580
rect 3152 31578 3176 31580
rect 3232 31578 3256 31580
rect 3312 31578 3318 31580
rect 3072 31526 3074 31578
rect 3254 31526 3256 31578
rect 3010 31524 3016 31526
rect 3072 31524 3096 31526
rect 3152 31524 3176 31526
rect 3232 31524 3256 31526
rect 3312 31524 3318 31526
rect 3010 31515 3318 31524
rect 2350 31036 2658 31045
rect 2350 31034 2356 31036
rect 2412 31034 2436 31036
rect 2492 31034 2516 31036
rect 2572 31034 2596 31036
rect 2652 31034 2658 31036
rect 2412 30982 2414 31034
rect 2594 30982 2596 31034
rect 2350 30980 2356 30982
rect 2412 30980 2436 30982
rect 2492 30980 2516 30982
rect 2572 30980 2596 30982
rect 2652 30980 2658 30982
rect 2350 30971 2658 30980
rect 4816 30802 4844 32166
rect 6012 31890 6040 35866
rect 6196 35834 6224 36178
rect 6184 35828 6236 35834
rect 6184 35770 6236 35776
rect 6092 35624 6144 35630
rect 6092 35566 6144 35572
rect 6104 33454 6132 35566
rect 6184 35012 6236 35018
rect 6184 34954 6236 34960
rect 6196 33998 6224 34954
rect 6184 33992 6236 33998
rect 6184 33934 6236 33940
rect 6092 33448 6144 33454
rect 6092 33390 6144 33396
rect 6000 31884 6052 31890
rect 6000 31826 6052 31832
rect 4804 30796 4856 30802
rect 4804 30738 4856 30744
rect 3010 30492 3318 30501
rect 3010 30490 3016 30492
rect 3072 30490 3096 30492
rect 3152 30490 3176 30492
rect 3232 30490 3256 30492
rect 3312 30490 3318 30492
rect 3072 30438 3074 30490
rect 3254 30438 3256 30490
rect 3010 30436 3016 30438
rect 3072 30436 3096 30438
rect 3152 30436 3176 30438
rect 3232 30436 3256 30438
rect 3312 30436 3318 30438
rect 3010 30427 3318 30436
rect 2350 29948 2658 29957
rect 2350 29946 2356 29948
rect 2412 29946 2436 29948
rect 2492 29946 2516 29948
rect 2572 29946 2596 29948
rect 2652 29946 2658 29948
rect 2412 29894 2414 29946
rect 2594 29894 2596 29946
rect 2350 29892 2356 29894
rect 2412 29892 2436 29894
rect 2492 29892 2516 29894
rect 2572 29892 2596 29894
rect 2652 29892 2658 29894
rect 2350 29883 2658 29892
rect 3010 29404 3318 29413
rect 3010 29402 3016 29404
rect 3072 29402 3096 29404
rect 3152 29402 3176 29404
rect 3232 29402 3256 29404
rect 3312 29402 3318 29404
rect 3072 29350 3074 29402
rect 3254 29350 3256 29402
rect 3010 29348 3016 29350
rect 3072 29348 3096 29350
rect 3152 29348 3176 29350
rect 3232 29348 3256 29350
rect 3312 29348 3318 29350
rect 3010 29339 3318 29348
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 2350 28860 2658 28869
rect 2350 28858 2356 28860
rect 2412 28858 2436 28860
rect 2492 28858 2516 28860
rect 2572 28858 2596 28860
rect 2652 28858 2658 28860
rect 2412 28806 2414 28858
rect 2594 28806 2596 28858
rect 2350 28804 2356 28806
rect 2412 28804 2436 28806
rect 2492 28804 2516 28806
rect 2572 28804 2596 28806
rect 2652 28804 2658 28806
rect 2350 28795 2658 28804
rect 3010 28316 3318 28325
rect 3010 28314 3016 28316
rect 3072 28314 3096 28316
rect 3152 28314 3176 28316
rect 3232 28314 3256 28316
rect 3312 28314 3318 28316
rect 3072 28262 3074 28314
rect 3254 28262 3256 28314
rect 3010 28260 3016 28262
rect 3072 28260 3096 28262
rect 3152 28260 3176 28262
rect 3232 28260 3256 28262
rect 3312 28260 3318 28262
rect 3010 28251 3318 28260
rect 4436 28076 4488 28082
rect 4436 28018 4488 28024
rect 2350 27772 2658 27781
rect 2350 27770 2356 27772
rect 2412 27770 2436 27772
rect 2492 27770 2516 27772
rect 2572 27770 2596 27772
rect 2652 27770 2658 27772
rect 2412 27718 2414 27770
rect 2594 27718 2596 27770
rect 2350 27716 2356 27718
rect 2412 27716 2436 27718
rect 2492 27716 2516 27718
rect 2572 27716 2596 27718
rect 2652 27716 2658 27718
rect 2350 27707 2658 27716
rect 3010 27228 3318 27237
rect 3010 27226 3016 27228
rect 3072 27226 3096 27228
rect 3152 27226 3176 27228
rect 3232 27226 3256 27228
rect 3312 27226 3318 27228
rect 3072 27174 3074 27226
rect 3254 27174 3256 27226
rect 3010 27172 3016 27174
rect 3072 27172 3096 27174
rect 3152 27172 3176 27174
rect 3232 27172 3256 27174
rect 3312 27172 3318 27174
rect 3010 27163 3318 27172
rect 2350 26684 2658 26693
rect 2350 26682 2356 26684
rect 2412 26682 2436 26684
rect 2492 26682 2516 26684
rect 2572 26682 2596 26684
rect 2652 26682 2658 26684
rect 2412 26630 2414 26682
rect 2594 26630 2596 26682
rect 2350 26628 2356 26630
rect 2412 26628 2436 26630
rect 2492 26628 2516 26630
rect 2572 26628 2596 26630
rect 2652 26628 2658 26630
rect 2350 26619 2658 26628
rect 4448 26450 4476 28018
rect 4724 28014 4752 28902
rect 4816 28626 4844 30738
rect 5080 30660 5132 30666
rect 5080 30602 5132 30608
rect 5092 30394 5120 30602
rect 5080 30388 5132 30394
rect 5080 30330 5132 30336
rect 5264 29504 5316 29510
rect 5264 29446 5316 29452
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5276 29306 5304 29446
rect 5264 29300 5316 29306
rect 5264 29242 5316 29248
rect 5920 29170 5948 29446
rect 5908 29164 5960 29170
rect 5908 29106 5960 29112
rect 5172 28960 5224 28966
rect 5172 28902 5224 28908
rect 5184 28626 5212 28902
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 5172 28620 5224 28626
rect 5172 28562 5224 28568
rect 4816 28218 4844 28562
rect 4804 28212 4856 28218
rect 4804 28154 4856 28160
rect 4712 28008 4764 28014
rect 4712 27950 4764 27956
rect 5724 26920 5776 26926
rect 5724 26862 5776 26868
rect 5736 26586 5764 26862
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 4436 26444 4488 26450
rect 4436 26386 4488 26392
rect 3010 26140 3318 26149
rect 3010 26138 3016 26140
rect 3072 26138 3096 26140
rect 3152 26138 3176 26140
rect 3232 26138 3256 26140
rect 3312 26138 3318 26140
rect 3072 26086 3074 26138
rect 3254 26086 3256 26138
rect 3010 26084 3016 26086
rect 3072 26084 3096 26086
rect 3152 26084 3176 26086
rect 3232 26084 3256 26086
rect 3312 26084 3318 26086
rect 3010 26075 3318 26084
rect 2350 25596 2658 25605
rect 2350 25594 2356 25596
rect 2412 25594 2436 25596
rect 2492 25594 2516 25596
rect 2572 25594 2596 25596
rect 2652 25594 2658 25596
rect 2412 25542 2414 25594
rect 2594 25542 2596 25594
rect 2350 25540 2356 25542
rect 2412 25540 2436 25542
rect 2492 25540 2516 25542
rect 2572 25540 2596 25542
rect 2652 25540 2658 25542
rect 2350 25531 2658 25540
rect 3010 25052 3318 25061
rect 3010 25050 3016 25052
rect 3072 25050 3096 25052
rect 3152 25050 3176 25052
rect 3232 25050 3256 25052
rect 3312 25050 3318 25052
rect 3072 24998 3074 25050
rect 3254 24998 3256 25050
rect 3010 24996 3016 24998
rect 3072 24996 3096 24998
rect 3152 24996 3176 24998
rect 3232 24996 3256 24998
rect 3312 24996 3318 24998
rect 3010 24987 3318 24996
rect 2350 24508 2658 24517
rect 2350 24506 2356 24508
rect 2412 24506 2436 24508
rect 2492 24506 2516 24508
rect 2572 24506 2596 24508
rect 2652 24506 2658 24508
rect 2412 24454 2414 24506
rect 2594 24454 2596 24506
rect 2350 24452 2356 24454
rect 2412 24452 2436 24454
rect 2492 24452 2516 24454
rect 2572 24452 2596 24454
rect 2652 24452 2658 24454
rect 2350 24443 2658 24452
rect 6012 24206 6040 31826
rect 6104 30326 6132 33390
rect 6184 32224 6236 32230
rect 6184 32166 6236 32172
rect 6196 31686 6224 32166
rect 6184 31680 6236 31686
rect 6184 31622 6236 31628
rect 6196 30394 6224 31622
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6092 30320 6144 30326
rect 6092 30262 6144 30268
rect 6104 29714 6132 30262
rect 6288 29714 6316 38966
rect 6564 38282 6592 39306
rect 6552 38276 6604 38282
rect 6552 38218 6604 38224
rect 6460 37868 6512 37874
rect 6460 37810 6512 37816
rect 6472 37466 6500 37810
rect 6460 37460 6512 37466
rect 6460 37402 6512 37408
rect 6460 36780 6512 36786
rect 6460 36722 6512 36728
rect 6472 36378 6500 36722
rect 6460 36372 6512 36378
rect 6460 36314 6512 36320
rect 6564 35894 6592 38218
rect 6748 37806 6776 39374
rect 6736 37800 6788 37806
rect 6736 37742 6788 37748
rect 6748 36718 6776 37742
rect 6736 36712 6788 36718
rect 6736 36654 6788 36660
rect 6564 35866 6684 35894
rect 6460 35080 6512 35086
rect 6460 35022 6512 35028
rect 6472 33658 6500 35022
rect 6552 33856 6604 33862
rect 6552 33798 6604 33804
rect 6460 33652 6512 33658
rect 6460 33594 6512 33600
rect 6564 33590 6592 33798
rect 6552 33584 6604 33590
rect 6552 33526 6604 33532
rect 6656 33402 6684 35866
rect 6748 35086 6776 36654
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 6748 34542 6776 35022
rect 6840 34610 6868 40326
rect 7024 40310 7236 40338
rect 7024 35894 7052 40310
rect 7760 39982 7788 41414
rect 7748 39976 7800 39982
rect 7748 39918 7800 39924
rect 7350 39740 7658 39749
rect 7350 39738 7356 39740
rect 7412 39738 7436 39740
rect 7492 39738 7516 39740
rect 7572 39738 7596 39740
rect 7652 39738 7658 39740
rect 7412 39686 7414 39738
rect 7594 39686 7596 39738
rect 7350 39684 7356 39686
rect 7412 39684 7436 39686
rect 7492 39684 7516 39686
rect 7572 39684 7596 39686
rect 7652 39684 7658 39686
rect 7350 39675 7658 39684
rect 7104 39364 7156 39370
rect 7104 39306 7156 39312
rect 7116 38418 7144 39306
rect 7656 39296 7708 39302
rect 7656 39238 7708 39244
rect 7668 39098 7696 39238
rect 7656 39092 7708 39098
rect 7656 39034 7708 39040
rect 7760 38826 7788 39918
rect 7196 38820 7248 38826
rect 7196 38762 7248 38768
rect 7748 38820 7800 38826
rect 7748 38762 7800 38768
rect 7104 38412 7156 38418
rect 7104 38354 7156 38360
rect 7104 37664 7156 37670
rect 7104 37606 7156 37612
rect 7116 37262 7144 37606
rect 7208 37330 7236 38762
rect 7350 38652 7658 38661
rect 7350 38650 7356 38652
rect 7412 38650 7436 38652
rect 7492 38650 7516 38652
rect 7572 38650 7596 38652
rect 7652 38650 7658 38652
rect 7412 38598 7414 38650
rect 7594 38598 7596 38650
rect 7350 38596 7356 38598
rect 7412 38596 7436 38598
rect 7492 38596 7516 38598
rect 7572 38596 7596 38598
rect 7652 38596 7658 38598
rect 7350 38587 7658 38596
rect 7748 38344 7800 38350
rect 7748 38286 7800 38292
rect 7760 37670 7788 38286
rect 7748 37664 7800 37670
rect 7748 37606 7800 37612
rect 7350 37564 7658 37573
rect 7350 37562 7356 37564
rect 7412 37562 7436 37564
rect 7492 37562 7516 37564
rect 7572 37562 7596 37564
rect 7652 37562 7658 37564
rect 7412 37510 7414 37562
rect 7594 37510 7596 37562
rect 7350 37508 7356 37510
rect 7412 37508 7436 37510
rect 7492 37508 7516 37510
rect 7572 37508 7596 37510
rect 7652 37508 7658 37510
rect 7350 37499 7658 37508
rect 7196 37324 7248 37330
rect 7196 37266 7248 37272
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 7208 36242 7236 37266
rect 7748 36712 7800 36718
rect 7748 36654 7800 36660
rect 7350 36476 7658 36485
rect 7350 36474 7356 36476
rect 7412 36474 7436 36476
rect 7492 36474 7516 36476
rect 7572 36474 7596 36476
rect 7652 36474 7658 36476
rect 7412 36422 7414 36474
rect 7594 36422 7596 36474
rect 7350 36420 7356 36422
rect 7412 36420 7436 36422
rect 7492 36420 7516 36422
rect 7572 36420 7596 36422
rect 7652 36420 7658 36422
rect 7350 36411 7658 36420
rect 7196 36236 7248 36242
rect 7196 36178 7248 36184
rect 6932 35866 7052 35894
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 6748 33862 6776 34478
rect 6736 33856 6788 33862
rect 6736 33798 6788 33804
rect 6564 33374 6684 33402
rect 6564 32434 6592 33374
rect 6460 32428 6512 32434
rect 6460 32370 6512 32376
rect 6552 32428 6604 32434
rect 6552 32370 6604 32376
rect 6472 32026 6500 32370
rect 6460 32020 6512 32026
rect 6460 31962 6512 31968
rect 6460 31340 6512 31346
rect 6460 31282 6512 31288
rect 6472 30938 6500 31282
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6460 30796 6512 30802
rect 6460 30738 6512 30744
rect 6472 30394 6500 30738
rect 6564 30734 6592 32370
rect 6748 32366 6776 33798
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6748 31278 6776 32302
rect 6736 31272 6788 31278
rect 6736 31214 6788 31220
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6460 30388 6512 30394
rect 6460 30330 6512 30336
rect 6092 29708 6144 29714
rect 6092 29650 6144 29656
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 6104 29102 6132 29650
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6104 28642 6132 29038
rect 6104 28614 6224 28642
rect 6092 28552 6144 28558
rect 6092 28494 6144 28500
rect 6104 28218 6132 28494
rect 6092 28212 6144 28218
rect 6092 28154 6144 28160
rect 6196 26926 6224 28614
rect 6288 28218 6316 29650
rect 6460 29640 6512 29646
rect 6460 29582 6512 29588
rect 6472 29306 6500 29582
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 6564 29186 6592 30670
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 6656 30190 6684 30534
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6656 29238 6684 30126
rect 6748 29646 6776 31214
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6472 29158 6592 29186
rect 6644 29232 6696 29238
rect 6644 29174 6696 29180
rect 6276 28212 6328 28218
rect 6276 28154 6328 28160
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6196 26466 6224 26862
rect 6368 26784 6420 26790
rect 6368 26726 6420 26732
rect 6104 26438 6224 26466
rect 6104 26042 6132 26438
rect 6184 26308 6236 26314
rect 6184 26250 6236 26256
rect 6196 26042 6224 26250
rect 6092 26036 6144 26042
rect 6092 25978 6144 25984
rect 6184 26036 6236 26042
rect 6184 25978 6236 25984
rect 6380 25770 6408 26726
rect 6368 25764 6420 25770
rect 6368 25706 6420 25712
rect 6000 24200 6052 24206
rect 6000 24142 6052 24148
rect 3010 23964 3318 23973
rect 3010 23962 3016 23964
rect 3072 23962 3096 23964
rect 3152 23962 3176 23964
rect 3232 23962 3256 23964
rect 3312 23962 3318 23964
rect 3072 23910 3074 23962
rect 3254 23910 3256 23962
rect 3010 23908 3016 23910
rect 3072 23908 3096 23910
rect 3152 23908 3176 23910
rect 3232 23908 3256 23910
rect 3312 23908 3318 23910
rect 3010 23899 3318 23908
rect 6472 23594 6500 29158
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6564 28422 6592 29038
rect 6748 28558 6776 29582
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6552 28416 6604 28422
rect 6552 28358 6604 28364
rect 6564 28150 6592 28358
rect 6552 28144 6604 28150
rect 6552 28086 6604 28092
rect 6748 26450 6776 28494
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6748 25702 6776 26386
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6736 25696 6788 25702
rect 6736 25638 6788 25644
rect 6656 25498 6684 25638
rect 6644 25492 6696 25498
rect 6644 25434 6696 25440
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6656 24614 6684 25094
rect 6748 24954 6776 25638
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6748 23610 6776 24142
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6656 23582 6776 23610
rect 2350 23420 2658 23429
rect 2350 23418 2356 23420
rect 2412 23418 2436 23420
rect 2492 23418 2516 23420
rect 2572 23418 2596 23420
rect 2652 23418 2658 23420
rect 2412 23366 2414 23418
rect 2594 23366 2596 23418
rect 2350 23364 2356 23366
rect 2412 23364 2436 23366
rect 2492 23364 2516 23366
rect 2572 23364 2596 23366
rect 2652 23364 2658 23366
rect 2350 23355 2658 23364
rect 3010 22876 3318 22885
rect 3010 22874 3016 22876
rect 3072 22874 3096 22876
rect 3152 22874 3176 22876
rect 3232 22874 3256 22876
rect 3312 22874 3318 22876
rect 3072 22822 3074 22874
rect 3254 22822 3256 22874
rect 3010 22820 3016 22822
rect 3072 22820 3096 22822
rect 3152 22820 3176 22822
rect 3232 22820 3256 22822
rect 3312 22820 3318 22822
rect 3010 22811 3318 22820
rect 2350 22332 2658 22341
rect 2350 22330 2356 22332
rect 2412 22330 2436 22332
rect 2492 22330 2516 22332
rect 2572 22330 2596 22332
rect 2652 22330 2658 22332
rect 2412 22278 2414 22330
rect 2594 22278 2596 22330
rect 2350 22276 2356 22278
rect 2412 22276 2436 22278
rect 2492 22276 2516 22278
rect 2572 22276 2596 22278
rect 2652 22276 2658 22278
rect 2350 22267 2658 22276
rect 3010 21788 3318 21797
rect 3010 21786 3016 21788
rect 3072 21786 3096 21788
rect 3152 21786 3176 21788
rect 3232 21786 3256 21788
rect 3312 21786 3318 21788
rect 3072 21734 3074 21786
rect 3254 21734 3256 21786
rect 3010 21732 3016 21734
rect 3072 21732 3096 21734
rect 3152 21732 3176 21734
rect 3232 21732 3256 21734
rect 3312 21732 3318 21734
rect 3010 21723 3318 21732
rect 2350 21244 2658 21253
rect 2350 21242 2356 21244
rect 2412 21242 2436 21244
rect 2492 21242 2516 21244
rect 2572 21242 2596 21244
rect 2652 21242 2658 21244
rect 2412 21190 2414 21242
rect 2594 21190 2596 21242
rect 2350 21188 2356 21190
rect 2412 21188 2436 21190
rect 2492 21188 2516 21190
rect 2572 21188 2596 21190
rect 2652 21188 2658 21190
rect 2350 21179 2658 21188
rect 3010 20700 3318 20709
rect 3010 20698 3016 20700
rect 3072 20698 3096 20700
rect 3152 20698 3176 20700
rect 3232 20698 3256 20700
rect 3312 20698 3318 20700
rect 3072 20646 3074 20698
rect 3254 20646 3256 20698
rect 3010 20644 3016 20646
rect 3072 20644 3096 20646
rect 3152 20644 3176 20646
rect 3232 20644 3256 20646
rect 3312 20644 3318 20646
rect 3010 20635 3318 20644
rect 2350 20156 2658 20165
rect 2350 20154 2356 20156
rect 2412 20154 2436 20156
rect 2492 20154 2516 20156
rect 2572 20154 2596 20156
rect 2652 20154 2658 20156
rect 2412 20102 2414 20154
rect 2594 20102 2596 20154
rect 2350 20100 2356 20102
rect 2412 20100 2436 20102
rect 2492 20100 2516 20102
rect 2572 20100 2596 20102
rect 2652 20100 2658 20102
rect 2350 20091 2658 20100
rect 3010 19612 3318 19621
rect 3010 19610 3016 19612
rect 3072 19610 3096 19612
rect 3152 19610 3176 19612
rect 3232 19610 3256 19612
rect 3312 19610 3318 19612
rect 3072 19558 3074 19610
rect 3254 19558 3256 19610
rect 3010 19556 3016 19558
rect 3072 19556 3096 19558
rect 3152 19556 3176 19558
rect 3232 19556 3256 19558
rect 3312 19556 3318 19558
rect 3010 19547 3318 19556
rect 2350 19068 2658 19077
rect 2350 19066 2356 19068
rect 2412 19066 2436 19068
rect 2492 19066 2516 19068
rect 2572 19066 2596 19068
rect 2652 19066 2658 19068
rect 2412 19014 2414 19066
rect 2594 19014 2596 19066
rect 2350 19012 2356 19014
rect 2412 19012 2436 19014
rect 2492 19012 2516 19014
rect 2572 19012 2596 19014
rect 2652 19012 2658 19014
rect 2350 19003 2658 19012
rect 3010 18524 3318 18533
rect 3010 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3176 18524
rect 3232 18522 3256 18524
rect 3312 18522 3318 18524
rect 3072 18470 3074 18522
rect 3254 18470 3256 18522
rect 3010 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3176 18470
rect 3232 18468 3256 18470
rect 3312 18468 3318 18470
rect 3010 18459 3318 18468
rect 2350 17980 2658 17989
rect 2350 17978 2356 17980
rect 2412 17978 2436 17980
rect 2492 17978 2516 17980
rect 2572 17978 2596 17980
rect 2652 17978 2658 17980
rect 2412 17926 2414 17978
rect 2594 17926 2596 17978
rect 2350 17924 2356 17926
rect 2412 17924 2436 17926
rect 2492 17924 2516 17926
rect 2572 17924 2596 17926
rect 2652 17924 2658 17926
rect 2350 17915 2658 17924
rect 3010 17436 3318 17445
rect 3010 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3176 17436
rect 3232 17434 3256 17436
rect 3312 17434 3318 17436
rect 3072 17382 3074 17434
rect 3254 17382 3256 17434
rect 3010 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3176 17382
rect 3232 17380 3256 17382
rect 3312 17380 3318 17382
rect 3010 17371 3318 17380
rect 2350 16892 2658 16901
rect 2350 16890 2356 16892
rect 2412 16890 2436 16892
rect 2492 16890 2516 16892
rect 2572 16890 2596 16892
rect 2652 16890 2658 16892
rect 2412 16838 2414 16890
rect 2594 16838 2596 16890
rect 2350 16836 2356 16838
rect 2412 16836 2436 16838
rect 2492 16836 2516 16838
rect 2572 16836 2596 16838
rect 2652 16836 2658 16838
rect 2350 16827 2658 16836
rect 3010 16348 3318 16357
rect 3010 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3176 16348
rect 3232 16346 3256 16348
rect 3312 16346 3318 16348
rect 3072 16294 3074 16346
rect 3254 16294 3256 16346
rect 3010 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3176 16294
rect 3232 16292 3256 16294
rect 3312 16292 3318 16294
rect 3010 16283 3318 16292
rect 2350 15804 2658 15813
rect 2350 15802 2356 15804
rect 2412 15802 2436 15804
rect 2492 15802 2516 15804
rect 2572 15802 2596 15804
rect 2652 15802 2658 15804
rect 2412 15750 2414 15802
rect 2594 15750 2596 15802
rect 2350 15748 2356 15750
rect 2412 15748 2436 15750
rect 2492 15748 2516 15750
rect 2572 15748 2596 15750
rect 2652 15748 2658 15750
rect 2350 15739 2658 15748
rect 3010 15260 3318 15269
rect 3010 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3176 15260
rect 3232 15258 3256 15260
rect 3312 15258 3318 15260
rect 3072 15206 3074 15258
rect 3254 15206 3256 15258
rect 3010 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3176 15206
rect 3232 15204 3256 15206
rect 3312 15204 3318 15206
rect 3010 15195 3318 15204
rect 2350 14716 2658 14725
rect 2350 14714 2356 14716
rect 2412 14714 2436 14716
rect 2492 14714 2516 14716
rect 2572 14714 2596 14716
rect 2652 14714 2658 14716
rect 2412 14662 2414 14714
rect 2594 14662 2596 14714
rect 2350 14660 2356 14662
rect 2412 14660 2436 14662
rect 2492 14660 2516 14662
rect 2572 14660 2596 14662
rect 2652 14660 2658 14662
rect 2350 14651 2658 14660
rect 6472 14346 6500 23530
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6564 22098 6592 23054
rect 6656 22438 6684 23582
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6748 23050 6776 23462
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6552 22092 6604 22098
rect 6552 22034 6604 22040
rect 6564 21010 6592 22034
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6564 19378 6592 20946
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6748 19446 6776 19926
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6564 18290 6592 19314
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6564 16658 6592 18226
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6656 16794 6684 17002
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6564 15162 6592 16594
rect 6748 16153 6776 17070
rect 6734 16144 6790 16153
rect 6734 16079 6790 16088
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 3010 14172 3318 14181
rect 3010 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3176 14172
rect 3232 14170 3256 14172
rect 3312 14170 3318 14172
rect 3072 14118 3074 14170
rect 3254 14118 3256 14170
rect 3010 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3176 14118
rect 3232 14116 3256 14118
rect 3312 14116 3318 14118
rect 3010 14107 3318 14116
rect 2350 13628 2658 13637
rect 2350 13626 2356 13628
rect 2412 13626 2436 13628
rect 2492 13626 2516 13628
rect 2572 13626 2596 13628
rect 2652 13626 2658 13628
rect 2412 13574 2414 13626
rect 2594 13574 2596 13626
rect 2350 13572 2356 13574
rect 2412 13572 2436 13574
rect 2492 13572 2516 13574
rect 2572 13572 2596 13574
rect 2652 13572 2658 13574
rect 2350 13563 2658 13572
rect 3010 13084 3318 13093
rect 3010 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3176 13084
rect 3232 13082 3256 13084
rect 3312 13082 3318 13084
rect 3072 13030 3074 13082
rect 3254 13030 3256 13082
rect 3010 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3176 13030
rect 3232 13028 3256 13030
rect 3312 13028 3318 13030
rect 3010 13019 3318 13028
rect 6104 12850 6132 14282
rect 6564 13938 6592 15098
rect 6656 15026 6684 15302
rect 6840 15094 6868 34546
rect 6932 31822 6960 35866
rect 7208 35034 7236 36178
rect 7350 35388 7658 35397
rect 7350 35386 7356 35388
rect 7412 35386 7436 35388
rect 7492 35386 7516 35388
rect 7572 35386 7596 35388
rect 7652 35386 7658 35388
rect 7412 35334 7414 35386
rect 7594 35334 7596 35386
rect 7350 35332 7356 35334
rect 7412 35332 7436 35334
rect 7492 35332 7516 35334
rect 7572 35332 7596 35334
rect 7652 35332 7658 35334
rect 7350 35323 7658 35332
rect 7760 35034 7788 36654
rect 7024 35006 7236 35034
rect 7300 35018 7788 35034
rect 7288 35012 7788 35018
rect 7024 34066 7052 35006
rect 7340 35006 7788 35012
rect 7288 34954 7340 34960
rect 7104 34944 7156 34950
rect 7300 34898 7328 34954
rect 7104 34886 7156 34892
rect 7012 34060 7064 34066
rect 7012 34002 7064 34008
rect 7012 33924 7064 33930
rect 7012 33866 7064 33872
rect 7024 33114 7052 33866
rect 7116 33658 7144 34886
rect 7208 34870 7328 34898
rect 7208 33862 7236 34870
rect 7350 34300 7658 34309
rect 7350 34298 7356 34300
rect 7412 34298 7436 34300
rect 7492 34298 7516 34300
rect 7572 34298 7596 34300
rect 7652 34298 7658 34300
rect 7412 34246 7414 34298
rect 7594 34246 7596 34298
rect 7350 34244 7356 34246
rect 7412 34244 7436 34246
rect 7492 34244 7516 34246
rect 7572 34244 7596 34246
rect 7652 34244 7658 34246
rect 7350 34235 7658 34244
rect 7380 34060 7432 34066
rect 7380 34002 7432 34008
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 7208 33538 7236 33798
rect 7116 33510 7236 33538
rect 7012 33108 7064 33114
rect 7012 33050 7064 33056
rect 7116 32502 7144 33510
rect 7392 33454 7420 34002
rect 7746 33552 7802 33561
rect 7746 33487 7802 33496
rect 7380 33448 7432 33454
rect 7380 33390 7432 33396
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 7208 32910 7236 33254
rect 7350 33212 7658 33221
rect 7350 33210 7356 33212
rect 7412 33210 7436 33212
rect 7492 33210 7516 33212
rect 7572 33210 7596 33212
rect 7652 33210 7658 33212
rect 7412 33158 7414 33210
rect 7594 33158 7596 33210
rect 7350 33156 7356 33158
rect 7412 33156 7436 33158
rect 7492 33156 7516 33158
rect 7572 33156 7596 33158
rect 7652 33156 7658 33158
rect 7350 33147 7658 33156
rect 7760 33114 7788 33487
rect 7748 33108 7800 33114
rect 7748 33050 7800 33056
rect 7196 32904 7248 32910
rect 7196 32846 7248 32852
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 7760 32230 7788 32778
rect 7104 32224 7156 32230
rect 7104 32166 7156 32172
rect 7748 32224 7800 32230
rect 7748 32166 7800 32172
rect 7116 31822 7144 32166
rect 7350 32124 7658 32133
rect 7350 32122 7356 32124
rect 7412 32122 7436 32124
rect 7492 32122 7516 32124
rect 7572 32122 7596 32124
rect 7652 32122 7658 32124
rect 7412 32070 7414 32122
rect 7594 32070 7596 32122
rect 7350 32068 7356 32070
rect 7412 32068 7436 32070
rect 7492 32068 7516 32070
rect 7572 32068 7596 32070
rect 7652 32068 7658 32070
rect 7350 32059 7658 32068
rect 7748 31884 7800 31890
rect 7748 31826 7800 31832
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7350 31036 7658 31045
rect 7350 31034 7356 31036
rect 7412 31034 7436 31036
rect 7492 31034 7516 31036
rect 7572 31034 7596 31036
rect 7652 31034 7658 31036
rect 7412 30982 7414 31034
rect 7594 30982 7596 31034
rect 7350 30980 7356 30982
rect 7412 30980 7436 30982
rect 7492 30980 7516 30982
rect 7572 30980 7596 30982
rect 7652 30980 7658 30982
rect 7350 30971 7658 30980
rect 7760 30802 7788 31826
rect 7748 30796 7800 30802
rect 7748 30738 7800 30744
rect 7350 29948 7658 29957
rect 7350 29946 7356 29948
rect 7412 29946 7436 29948
rect 7492 29946 7516 29948
rect 7572 29946 7596 29948
rect 7652 29946 7658 29948
rect 7412 29894 7414 29946
rect 7594 29894 7596 29946
rect 7350 29892 7356 29894
rect 7412 29892 7436 29894
rect 7492 29892 7516 29894
rect 7572 29892 7596 29894
rect 7652 29892 7658 29894
rect 7350 29883 7658 29892
rect 7760 29102 7788 30738
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 7012 28484 7064 28490
rect 7012 28426 7064 28432
rect 7024 28218 7052 28426
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7116 28098 7144 28562
rect 7024 28070 7144 28098
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6932 26586 6960 26862
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 7024 26466 7052 28070
rect 7208 28014 7236 28970
rect 7350 28860 7658 28869
rect 7350 28858 7356 28860
rect 7412 28858 7436 28860
rect 7492 28858 7516 28860
rect 7572 28858 7596 28860
rect 7652 28858 7658 28860
rect 7412 28806 7414 28858
rect 7594 28806 7596 28858
rect 7350 28804 7356 28806
rect 7412 28804 7436 28806
rect 7492 28804 7516 28806
rect 7572 28804 7596 28806
rect 7652 28804 7658 28806
rect 7350 28795 7658 28804
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7350 27772 7658 27781
rect 7350 27770 7356 27772
rect 7412 27770 7436 27772
rect 7492 27770 7516 27772
rect 7572 27770 7596 27772
rect 7652 27770 7658 27772
rect 7412 27718 7414 27770
rect 7594 27718 7596 27770
rect 7350 27716 7356 27718
rect 7412 27716 7436 27718
rect 7492 27716 7516 27718
rect 7572 27716 7596 27718
rect 7652 27716 7658 27718
rect 7350 27707 7658 27716
rect 7852 27418 7880 41482
rect 8010 41372 8318 41381
rect 8010 41370 8016 41372
rect 8072 41370 8096 41372
rect 8152 41370 8176 41372
rect 8232 41370 8256 41372
rect 8312 41370 8318 41372
rect 8072 41318 8074 41370
rect 8254 41318 8256 41370
rect 8010 41316 8016 41318
rect 8072 41316 8096 41318
rect 8152 41316 8176 41318
rect 8232 41316 8256 41318
rect 8312 41316 8318 41318
rect 8010 41307 8318 41316
rect 8392 40928 8444 40934
rect 8392 40870 8444 40876
rect 8404 40633 8432 40870
rect 8390 40624 8446 40633
rect 8390 40559 8446 40568
rect 8010 40284 8318 40293
rect 8010 40282 8016 40284
rect 8072 40282 8096 40284
rect 8152 40282 8176 40284
rect 8232 40282 8256 40284
rect 8312 40282 8318 40284
rect 8072 40230 8074 40282
rect 8254 40230 8256 40282
rect 8010 40228 8016 40230
rect 8072 40228 8096 40230
rect 8152 40228 8176 40230
rect 8232 40228 8256 40230
rect 8312 40228 8318 40230
rect 8010 40219 8318 40228
rect 8390 39264 8446 39273
rect 8010 39196 8318 39205
rect 8390 39199 8446 39208
rect 8010 39194 8016 39196
rect 8072 39194 8096 39196
rect 8152 39194 8176 39196
rect 8232 39194 8256 39196
rect 8312 39194 8318 39196
rect 8072 39142 8074 39194
rect 8254 39142 8256 39194
rect 8010 39140 8016 39142
rect 8072 39140 8096 39142
rect 8152 39140 8176 39142
rect 8232 39140 8256 39142
rect 8312 39140 8318 39142
rect 8010 39131 8318 39140
rect 8404 39098 8432 39199
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8392 38208 8444 38214
rect 8392 38150 8444 38156
rect 8010 38108 8318 38117
rect 8010 38106 8016 38108
rect 8072 38106 8096 38108
rect 8152 38106 8176 38108
rect 8232 38106 8256 38108
rect 8312 38106 8318 38108
rect 8072 38054 8074 38106
rect 8254 38054 8256 38106
rect 8010 38052 8016 38054
rect 8072 38052 8096 38054
rect 8152 38052 8176 38054
rect 8232 38052 8256 38054
rect 8312 38052 8318 38054
rect 8010 38043 8318 38052
rect 8024 37936 8076 37942
rect 8404 37913 8432 38150
rect 8024 37878 8076 37884
rect 8390 37904 8446 37913
rect 8036 37210 8064 37878
rect 8390 37839 8446 37848
rect 7944 37182 8064 37210
rect 7944 36922 7972 37182
rect 8010 37020 8318 37029
rect 8010 37018 8016 37020
rect 8072 37018 8096 37020
rect 8152 37018 8176 37020
rect 8232 37018 8256 37020
rect 8312 37018 8318 37020
rect 8072 36966 8074 37018
rect 8254 36966 8256 37018
rect 8010 36964 8016 36966
rect 8072 36964 8096 36966
rect 8152 36964 8176 36966
rect 8232 36964 8256 36966
rect 8312 36964 8318 36966
rect 8010 36955 8318 36964
rect 7932 36916 7984 36922
rect 7932 36858 7984 36864
rect 8390 36544 8446 36553
rect 8390 36479 8446 36488
rect 8404 36378 8432 36479
rect 8392 36372 8444 36378
rect 8392 36314 8444 36320
rect 8010 35932 8318 35941
rect 8010 35930 8016 35932
rect 8072 35930 8096 35932
rect 8152 35930 8176 35932
rect 8232 35930 8256 35932
rect 8312 35930 8318 35932
rect 8072 35878 8074 35930
rect 8254 35878 8256 35930
rect 8010 35876 8016 35878
rect 8072 35876 8096 35878
rect 8152 35876 8176 35878
rect 8232 35876 8256 35878
rect 8312 35876 8318 35878
rect 8010 35867 8318 35876
rect 8024 35692 8076 35698
rect 8024 35634 8076 35640
rect 8036 34950 8064 35634
rect 8392 35488 8444 35494
rect 8392 35430 8444 35436
rect 8404 35193 8432 35430
rect 8390 35184 8446 35193
rect 8390 35119 8446 35128
rect 8024 34944 8076 34950
rect 8024 34886 8076 34892
rect 8010 34844 8318 34853
rect 8010 34842 8016 34844
rect 8072 34842 8096 34844
rect 8152 34842 8176 34844
rect 8232 34842 8256 34844
rect 8312 34842 8318 34844
rect 8072 34790 8074 34842
rect 8254 34790 8256 34842
rect 8010 34788 8016 34790
rect 8072 34788 8096 34790
rect 8152 34788 8176 34790
rect 8232 34788 8256 34790
rect 8312 34788 8318 34790
rect 8010 34779 8318 34788
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7944 33658 7972 33798
rect 8010 33756 8318 33765
rect 8010 33754 8016 33756
rect 8072 33754 8096 33756
rect 8152 33754 8176 33756
rect 8232 33754 8256 33756
rect 8312 33754 8318 33756
rect 8072 33702 8074 33754
rect 8254 33702 8256 33754
rect 8010 33700 8016 33702
rect 8072 33700 8096 33702
rect 8152 33700 8176 33702
rect 8232 33700 8256 33702
rect 8312 33700 8318 33702
rect 8010 33691 8318 33700
rect 7932 33652 7984 33658
rect 7932 33594 7984 33600
rect 7944 33114 7972 33594
rect 8024 33448 8076 33454
rect 8024 33390 8076 33396
rect 7932 33108 7984 33114
rect 7932 33050 7984 33056
rect 8036 32858 8064 33390
rect 7944 32830 8064 32858
rect 7944 31890 7972 32830
rect 8668 32768 8720 32774
rect 8668 32710 8720 32716
rect 8010 32668 8318 32677
rect 8010 32666 8016 32668
rect 8072 32666 8096 32668
rect 8152 32666 8176 32668
rect 8232 32666 8256 32668
rect 8312 32666 8318 32668
rect 8072 32614 8074 32666
rect 8254 32614 8256 32666
rect 8010 32612 8016 32614
rect 8072 32612 8096 32614
rect 8152 32612 8176 32614
rect 8232 32612 8256 32614
rect 8312 32612 8318 32614
rect 8010 32603 8318 32612
rect 8680 32473 8708 32710
rect 8666 32464 8722 32473
rect 8666 32399 8722 32408
rect 7932 31884 7984 31890
rect 7932 31826 7984 31832
rect 8010 31580 8318 31589
rect 8010 31578 8016 31580
rect 8072 31578 8096 31580
rect 8152 31578 8176 31580
rect 8232 31578 8256 31580
rect 8312 31578 8318 31580
rect 8072 31526 8074 31578
rect 8254 31526 8256 31578
rect 8010 31524 8016 31526
rect 8072 31524 8096 31526
rect 8152 31524 8176 31526
rect 8232 31524 8256 31526
rect 8312 31524 8318 31526
rect 8010 31515 8318 31524
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 8036 30938 8064 31350
rect 8390 31104 8446 31113
rect 8390 31039 8446 31048
rect 8404 30938 8432 31039
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 8392 30932 8444 30938
rect 8392 30874 8444 30880
rect 8036 30682 8064 30874
rect 7944 30654 8064 30682
rect 7944 29730 7972 30654
rect 8010 30492 8318 30501
rect 8010 30490 8016 30492
rect 8072 30490 8096 30492
rect 8152 30490 8176 30492
rect 8232 30490 8256 30492
rect 8312 30490 8318 30492
rect 8072 30438 8074 30490
rect 8254 30438 8256 30490
rect 8010 30436 8016 30438
rect 8072 30436 8096 30438
rect 8152 30436 8176 30438
rect 8232 30436 8256 30438
rect 8312 30436 8318 30438
rect 8010 30427 8318 30436
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 8404 29753 8432 29990
rect 8390 29744 8446 29753
rect 7944 29702 8064 29730
rect 7944 28642 7972 29702
rect 8036 29646 8064 29702
rect 8390 29679 8446 29688
rect 8024 29640 8076 29646
rect 8024 29582 8076 29588
rect 8010 29404 8318 29413
rect 8010 29402 8016 29404
rect 8072 29402 8096 29404
rect 8152 29402 8176 29404
rect 8232 29402 8256 29404
rect 8312 29402 8318 29404
rect 8072 29350 8074 29402
rect 8254 29350 8256 29402
rect 8010 29348 8016 29350
rect 8072 29348 8096 29350
rect 8152 29348 8176 29350
rect 8232 29348 8256 29350
rect 8312 29348 8318 29350
rect 8010 29339 8318 29348
rect 7944 28614 8064 28642
rect 8036 28558 8064 28614
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 8390 28384 8446 28393
rect 8010 28316 8318 28325
rect 8390 28319 8446 28328
rect 8010 28314 8016 28316
rect 8072 28314 8096 28316
rect 8152 28314 8176 28316
rect 8232 28314 8256 28316
rect 8312 28314 8318 28316
rect 8072 28262 8074 28314
rect 8254 28262 8256 28314
rect 8010 28260 8016 28262
rect 8072 28260 8096 28262
rect 8152 28260 8176 28262
rect 8232 28260 8256 28262
rect 8312 28260 8318 28262
rect 8010 28251 8318 28260
rect 8404 28218 8432 28319
rect 8392 28212 8444 28218
rect 8392 28154 8444 28160
rect 6932 26450 7052 26466
rect 6920 26444 7052 26450
rect 6972 26438 7052 26444
rect 6920 26386 6972 26392
rect 7024 25906 7052 26438
rect 7116 27390 7880 27418
rect 7932 27396 7984 27402
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7024 24954 7052 25842
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7116 23746 7144 27390
rect 7932 27338 7984 27344
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7208 25498 7236 26930
rect 7350 26684 7658 26693
rect 7350 26682 7356 26684
rect 7412 26682 7436 26684
rect 7492 26682 7516 26684
rect 7572 26682 7596 26684
rect 7652 26682 7658 26684
rect 7412 26630 7414 26682
rect 7594 26630 7596 26682
rect 7350 26628 7356 26630
rect 7412 26628 7436 26630
rect 7492 26628 7516 26630
rect 7572 26628 7596 26630
rect 7652 26628 7658 26630
rect 7350 26619 7658 26628
rect 7760 26586 7788 26930
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7760 25673 7788 26318
rect 7746 25664 7802 25673
rect 7350 25596 7658 25605
rect 7746 25599 7802 25608
rect 7350 25594 7356 25596
rect 7412 25594 7436 25596
rect 7492 25594 7516 25596
rect 7572 25594 7596 25596
rect 7652 25594 7658 25596
rect 7412 25542 7414 25594
rect 7594 25542 7596 25594
rect 7350 25540 7356 25542
rect 7412 25540 7436 25542
rect 7492 25540 7516 25542
rect 7572 25540 7596 25542
rect 7652 25540 7658 25542
rect 7350 25531 7658 25540
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7208 24410 7236 25434
rect 7852 25362 7880 27270
rect 7944 27010 7972 27338
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8010 27228 8318 27237
rect 8010 27226 8016 27228
rect 8072 27226 8096 27228
rect 8152 27226 8176 27228
rect 8232 27226 8256 27228
rect 8312 27226 8318 27228
rect 8072 27174 8074 27226
rect 8254 27174 8256 27226
rect 8010 27172 8016 27174
rect 8072 27172 8096 27174
rect 8152 27172 8176 27174
rect 8232 27172 8256 27174
rect 8312 27172 8318 27174
rect 8010 27163 8318 27172
rect 8404 27130 8432 27270
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8864 27033 8892 27270
rect 8850 27024 8906 27033
rect 7944 26982 8064 27010
rect 7932 26784 7984 26790
rect 7932 26726 7984 26732
rect 7944 26042 7972 26726
rect 8036 26382 8064 26982
rect 8850 26959 8906 26968
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8010 26140 8318 26149
rect 8010 26138 8016 26140
rect 8072 26138 8096 26140
rect 8152 26138 8176 26140
rect 8232 26138 8256 26140
rect 8312 26138 8318 26140
rect 8072 26086 8074 26138
rect 8254 26086 8256 26138
rect 8010 26084 8016 26086
rect 8072 26084 8096 26086
rect 8152 26084 8176 26086
rect 8232 26084 8256 26086
rect 8312 26084 8318 26086
rect 8010 26075 8318 26084
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 7840 25356 7892 25362
rect 7840 25298 7892 25304
rect 8010 25052 8318 25061
rect 8010 25050 8016 25052
rect 8072 25050 8096 25052
rect 8152 25050 8176 25052
rect 8232 25050 8256 25052
rect 8312 25050 8318 25052
rect 8072 24998 8074 25050
rect 8254 24998 8256 25050
rect 8010 24996 8016 24998
rect 8072 24996 8096 24998
rect 8152 24996 8176 24998
rect 8232 24996 8256 24998
rect 8312 24996 8318 24998
rect 8010 24987 8318 24996
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 7350 24508 7658 24517
rect 7350 24506 7356 24508
rect 7412 24506 7436 24508
rect 7492 24506 7516 24508
rect 7572 24506 7596 24508
rect 7652 24506 7658 24508
rect 7412 24454 7414 24506
rect 7594 24454 7596 24506
rect 7350 24452 7356 24454
rect 7412 24452 7436 24454
rect 7492 24452 7516 24454
rect 7572 24452 7596 24454
rect 7652 24452 7658 24454
rect 7350 24443 7658 24452
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7378 24304 7434 24313
rect 7024 23718 7144 23746
rect 7208 24262 7378 24290
rect 6920 23044 6972 23050
rect 6920 22986 6972 22992
rect 6932 22030 6960 22986
rect 7024 22522 7052 23718
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7116 23050 7144 23530
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7208 22658 7236 24262
rect 7378 24239 7434 24248
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 7760 23866 7788 24006
rect 7852 23866 7880 24006
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7350 23420 7658 23429
rect 7350 23418 7356 23420
rect 7412 23418 7436 23420
rect 7492 23418 7516 23420
rect 7572 23418 7596 23420
rect 7652 23418 7658 23420
rect 7412 23366 7414 23418
rect 7594 23366 7596 23418
rect 7350 23364 7356 23366
rect 7412 23364 7436 23366
rect 7492 23364 7516 23366
rect 7572 23364 7596 23366
rect 7652 23364 7658 23366
rect 7350 23355 7658 23364
rect 7852 22778 7880 23462
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7380 22704 7432 22710
rect 7208 22642 7328 22658
rect 7380 22646 7432 22652
rect 7208 22636 7340 22642
rect 7208 22630 7288 22636
rect 7288 22578 7340 22584
rect 7392 22522 7420 22646
rect 7944 22624 7972 24074
rect 8010 23964 8318 23973
rect 8010 23962 8016 23964
rect 8072 23962 8096 23964
rect 8152 23962 8176 23964
rect 8232 23962 8256 23964
rect 8312 23962 8318 23964
rect 8072 23910 8074 23962
rect 8254 23910 8256 23962
rect 8010 23908 8016 23910
rect 8072 23908 8096 23910
rect 8152 23908 8176 23910
rect 8232 23908 8256 23910
rect 8312 23908 8318 23910
rect 8010 23899 8318 23908
rect 8404 23866 8432 24550
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8312 23322 8340 23598
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8390 22944 8446 22953
rect 8010 22876 8318 22885
rect 8390 22879 8446 22888
rect 8010 22874 8016 22876
rect 8072 22874 8096 22876
rect 8152 22874 8176 22876
rect 8232 22874 8256 22876
rect 8312 22874 8318 22876
rect 8072 22822 8074 22874
rect 8254 22822 8256 22874
rect 8010 22820 8016 22822
rect 8072 22820 8096 22822
rect 8152 22820 8176 22822
rect 8232 22820 8256 22822
rect 8312 22820 8318 22822
rect 8010 22811 8318 22820
rect 8404 22778 8432 22879
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 7024 22494 7144 22522
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7024 22094 7052 22374
rect 7116 22250 7144 22494
rect 7300 22494 7420 22522
rect 7852 22596 7972 22624
rect 7852 22506 7880 22596
rect 7840 22500 7892 22506
rect 7300 22438 7328 22494
rect 7840 22442 7892 22448
rect 7932 22500 7984 22506
rect 7932 22442 7984 22448
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7350 22332 7658 22341
rect 7350 22330 7356 22332
rect 7412 22330 7436 22332
rect 7492 22330 7516 22332
rect 7572 22330 7596 22332
rect 7652 22330 7658 22332
rect 7412 22278 7414 22330
rect 7594 22278 7596 22330
rect 7350 22276 7356 22278
rect 7412 22276 7436 22278
rect 7492 22276 7516 22278
rect 7572 22276 7596 22278
rect 7652 22276 7658 22278
rect 7350 22267 7658 22276
rect 7116 22222 7236 22250
rect 7024 22066 7144 22094
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 21146 6960 21966
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 7024 21554 7052 21830
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 7116 21026 7144 22066
rect 6932 20998 7144 21026
rect 6932 17610 6960 20998
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7116 20602 7144 20810
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7208 20482 7236 22222
rect 7760 21962 7788 22374
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7944 21486 7972 22442
rect 8010 21788 8318 21797
rect 8010 21786 8016 21788
rect 8072 21786 8096 21788
rect 8152 21786 8176 21788
rect 8232 21786 8256 21788
rect 8312 21786 8318 21788
rect 8072 21734 8074 21786
rect 8254 21734 8256 21786
rect 8010 21732 8016 21734
rect 8072 21732 8096 21734
rect 8152 21732 8176 21734
rect 8232 21732 8256 21734
rect 8312 21732 8318 21734
rect 8010 21723 8318 21732
rect 8300 21616 8352 21622
rect 8298 21584 8300 21593
rect 8352 21584 8354 21593
rect 8298 21519 8354 21528
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 7350 21244 7658 21253
rect 7350 21242 7356 21244
rect 7412 21242 7436 21244
rect 7492 21242 7516 21244
rect 7572 21242 7596 21244
rect 7652 21242 7658 21244
rect 7412 21190 7414 21242
rect 7594 21190 7596 21242
rect 7350 21188 7356 21190
rect 7412 21188 7436 21190
rect 7492 21188 7516 21190
rect 7572 21188 7596 21190
rect 7652 21188 7658 21190
rect 7350 21179 7658 21188
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7300 20874 7328 21082
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7024 20454 7236 20482
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 16114 6960 16934
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6840 14414 6868 15030
rect 6932 14618 6960 15438
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 14006 6960 14214
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 7024 13818 7052 20454
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7116 19530 7144 20198
rect 7208 19718 7236 20334
rect 7300 20262 7328 20810
rect 7760 20602 7788 21286
rect 7944 20602 7972 21422
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8010 20700 8318 20709
rect 8010 20698 8016 20700
rect 8072 20698 8096 20700
rect 8152 20698 8176 20700
rect 8232 20698 8256 20700
rect 8312 20698 8318 20700
rect 8072 20646 8074 20698
rect 8254 20646 8256 20698
rect 8010 20644 8016 20646
rect 8072 20644 8096 20646
rect 8152 20644 8176 20646
rect 8232 20644 8256 20646
rect 8312 20644 8318 20646
rect 8010 20635 8318 20644
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7350 20156 7658 20165
rect 7350 20154 7356 20156
rect 7412 20154 7436 20156
rect 7492 20154 7516 20156
rect 7572 20154 7596 20156
rect 7652 20154 7658 20156
rect 7412 20102 7414 20154
rect 7594 20102 7596 20154
rect 7350 20100 7356 20102
rect 7412 20100 7436 20102
rect 7492 20100 7516 20102
rect 7572 20100 7596 20102
rect 7652 20100 7658 20102
rect 7350 20091 7658 20100
rect 7760 20058 7788 20198
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7852 19802 7880 20266
rect 7760 19774 7880 19802
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7116 19514 7236 19530
rect 7116 19508 7248 19514
rect 7116 19502 7196 19508
rect 7196 19450 7248 19456
rect 7208 18850 7236 19450
rect 7350 19068 7658 19077
rect 7350 19066 7356 19068
rect 7412 19066 7436 19068
rect 7492 19066 7516 19068
rect 7572 19066 7596 19068
rect 7652 19066 7658 19068
rect 7412 19014 7414 19066
rect 7594 19014 7596 19066
rect 7350 19012 7356 19014
rect 7412 19012 7436 19014
rect 7492 19012 7516 19014
rect 7572 19012 7596 19014
rect 7652 19012 7658 19014
rect 7350 19003 7658 19012
rect 7208 18822 7328 18850
rect 7760 18834 7788 19774
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18426 7236 18566
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7300 18222 7328 18822
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7852 18766 7880 19654
rect 7944 19394 7972 20402
rect 8128 20058 8156 20402
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8220 19718 8248 20470
rect 8298 20224 8354 20233
rect 8298 20159 8354 20168
rect 8312 19786 8340 20159
rect 8404 19922 8432 20742
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8010 19612 8318 19621
rect 8010 19610 8016 19612
rect 8072 19610 8096 19612
rect 8152 19610 8176 19612
rect 8232 19610 8256 19612
rect 8312 19610 8318 19612
rect 8072 19558 8074 19610
rect 8254 19558 8256 19610
rect 8010 19556 8016 19558
rect 8072 19556 8096 19558
rect 8152 19556 8176 19558
rect 8232 19556 8256 19558
rect 8312 19556 8318 19558
rect 8010 19547 8318 19556
rect 8404 19394 8432 19654
rect 7944 19366 8064 19394
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 8036 18850 8064 19366
rect 8220 19366 8432 19394
rect 8220 18970 8248 19366
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8206 18864 8262 18873
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7944 18442 7972 18838
rect 8036 18822 8206 18850
rect 8206 18799 8262 18808
rect 8010 18524 8318 18533
rect 8010 18522 8016 18524
rect 8072 18522 8096 18524
rect 8152 18522 8176 18524
rect 8232 18522 8256 18524
rect 8312 18522 8318 18524
rect 8072 18470 8074 18522
rect 8254 18470 8256 18522
rect 8010 18468 8016 18470
rect 8072 18468 8096 18470
rect 8152 18468 8176 18470
rect 8232 18468 8256 18470
rect 8312 18468 8318 18470
rect 8010 18459 8318 18468
rect 7852 18414 7972 18442
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7350 17980 7658 17989
rect 7350 17978 7356 17980
rect 7412 17978 7436 17980
rect 7492 17978 7516 17980
rect 7572 17978 7596 17980
rect 7652 17978 7658 17980
rect 7412 17926 7414 17978
rect 7594 17926 7596 17978
rect 7350 17924 7356 17926
rect 7412 17924 7436 17926
rect 7492 17924 7516 17926
rect 7572 17924 7596 17926
rect 7652 17924 7658 17926
rect 7350 17915 7658 17924
rect 7852 17882 7880 18414
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 6932 13790 7052 13818
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12986 6776 13126
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 2350 12540 2658 12549
rect 2350 12538 2356 12540
rect 2412 12538 2436 12540
rect 2492 12538 2516 12540
rect 2572 12538 2596 12540
rect 2652 12538 2658 12540
rect 2412 12486 2414 12538
rect 2594 12486 2596 12538
rect 2350 12484 2356 12486
rect 2412 12484 2436 12486
rect 2492 12484 2516 12486
rect 2572 12484 2596 12486
rect 2652 12484 2658 12486
rect 2350 12475 2658 12484
rect 3010 11996 3318 12005
rect 3010 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3176 11996
rect 3232 11994 3256 11996
rect 3312 11994 3318 11996
rect 3072 11942 3074 11994
rect 3254 11942 3256 11994
rect 3010 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3176 11942
rect 3232 11940 3256 11942
rect 3312 11940 3318 11942
rect 3010 11931 3318 11940
rect 2350 11452 2658 11461
rect 2350 11450 2356 11452
rect 2412 11450 2436 11452
rect 2492 11450 2516 11452
rect 2572 11450 2596 11452
rect 2652 11450 2658 11452
rect 2412 11398 2414 11450
rect 2594 11398 2596 11450
rect 2350 11396 2356 11398
rect 2412 11396 2436 11398
rect 2492 11396 2516 11398
rect 2572 11396 2596 11398
rect 2652 11396 2658 11398
rect 2350 11387 2658 11396
rect 6564 11218 6592 12786
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 11898 6776 12106
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11218 6868 11494
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 3010 10908 3318 10917
rect 3010 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3176 10908
rect 3232 10906 3256 10908
rect 3312 10906 3318 10908
rect 3072 10854 3074 10906
rect 3254 10854 3256 10906
rect 3010 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3176 10854
rect 3232 10852 3256 10854
rect 3312 10852 3318 10854
rect 3010 10843 3318 10852
rect 2350 10364 2658 10373
rect 2350 10362 2356 10364
rect 2412 10362 2436 10364
rect 2492 10362 2516 10364
rect 2572 10362 2596 10364
rect 2652 10362 2658 10364
rect 2412 10310 2414 10362
rect 2594 10310 2596 10362
rect 2350 10308 2356 10310
rect 2412 10308 2436 10310
rect 2492 10308 2516 10310
rect 2572 10308 2596 10310
rect 2652 10308 2658 10310
rect 2350 10299 2658 10308
rect 6564 10130 6592 11154
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 3010 9820 3318 9829
rect 3010 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3176 9820
rect 3232 9818 3256 9820
rect 3312 9818 3318 9820
rect 3072 9766 3074 9818
rect 3254 9766 3256 9818
rect 3010 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3176 9766
rect 3232 9764 3256 9766
rect 3312 9764 3318 9766
rect 3010 9755 3318 9764
rect 2350 9276 2658 9285
rect 2350 9274 2356 9276
rect 2412 9274 2436 9276
rect 2492 9274 2516 9276
rect 2572 9274 2596 9276
rect 2652 9274 2658 9276
rect 2412 9222 2414 9274
rect 2594 9222 2596 9274
rect 2350 9220 2356 9222
rect 2412 9220 2436 9222
rect 2492 9220 2516 9222
rect 2572 9220 2596 9222
rect 2652 9220 2658 9222
rect 2350 9211 2658 9220
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 6564 8498 6592 10066
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6748 9178 6776 9454
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 2350 8188 2658 8197
rect 2350 8186 2356 8188
rect 2412 8186 2436 8188
rect 2492 8186 2516 8188
rect 2572 8186 2596 8188
rect 2652 8186 2658 8188
rect 2412 8134 2414 8186
rect 2594 8134 2596 8186
rect 2350 8132 2356 8134
rect 2412 8132 2436 8134
rect 2492 8132 2516 8134
rect 2572 8132 2596 8134
rect 2652 8132 2658 8134
rect 2350 8123 2658 8132
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 3988 7342 4016 7890
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4172 7546 4200 7754
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7546 4476 7686
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4816 7478 4844 7958
rect 5092 7886 5120 8230
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5368 7818 5672 7834
rect 5356 7812 5672 7818
rect 5408 7806 5672 7812
rect 5356 7754 5408 7760
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 2350 7100 2658 7109
rect 2350 7098 2356 7100
rect 2412 7098 2436 7100
rect 2492 7098 2516 7100
rect 2572 7098 2596 7100
rect 2652 7098 2658 7100
rect 2412 7046 2414 7098
rect 2594 7046 2596 7098
rect 2350 7044 2356 7046
rect 2412 7044 2436 7046
rect 2492 7044 2516 7046
rect 2572 7044 2596 7046
rect 2652 7044 2658 7046
rect 2350 7035 2658 7044
rect 3896 7002 3924 7142
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3988 6730 4016 7278
rect 4816 6730 4844 7414
rect 5552 7002 5580 7686
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6730 5672 7806
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7546 5764 7754
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 6012 7342 6040 8366
rect 6564 8022 6592 8434
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6564 7410 6592 7958
rect 6932 7818 6960 13790
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7024 11014 7052 12922
rect 7116 12866 7144 17478
rect 7760 17338 7788 17478
rect 7852 17338 7880 17478
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7944 17218 7972 18226
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8010 17436 8318 17445
rect 8010 17434 8016 17436
rect 8072 17434 8096 17436
rect 8152 17434 8176 17436
rect 8232 17434 8256 17436
rect 8312 17434 8318 17436
rect 8072 17382 8074 17434
rect 8254 17382 8256 17434
rect 8010 17380 8016 17382
rect 8072 17380 8096 17382
rect 8152 17380 8176 17382
rect 8232 17380 8256 17382
rect 8312 17380 8318 17382
rect 8010 17371 8318 17380
rect 7852 17190 7972 17218
rect 8404 17202 8432 18022
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8496 17513 8524 17546
rect 8482 17504 8538 17513
rect 8482 17439 8538 17448
rect 8392 17196 8444 17202
rect 7350 16892 7658 16901
rect 7350 16890 7356 16892
rect 7412 16890 7436 16892
rect 7492 16890 7516 16892
rect 7572 16890 7596 16892
rect 7652 16890 7658 16892
rect 7412 16838 7414 16890
rect 7594 16838 7596 16890
rect 7350 16836 7356 16838
rect 7412 16836 7436 16838
rect 7492 16836 7516 16838
rect 7572 16836 7596 16838
rect 7652 16836 7658 16838
rect 7350 16827 7658 16836
rect 7852 16522 7880 17190
rect 8392 17138 8444 17144
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7944 16250 7972 16934
rect 8312 16794 8340 17070
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8010 16348 8318 16357
rect 8010 16346 8016 16348
rect 8072 16346 8096 16348
rect 8152 16346 8176 16348
rect 8232 16346 8256 16348
rect 8312 16346 8318 16348
rect 8072 16294 8074 16346
rect 8254 16294 8256 16346
rect 8010 16292 8016 16294
rect 8072 16292 8096 16294
rect 8152 16292 8176 16294
rect 8232 16292 8256 16294
rect 8312 16292 8318 16294
rect 8010 16283 8318 16292
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7350 15804 7658 15813
rect 7350 15802 7356 15804
rect 7412 15802 7436 15804
rect 7492 15802 7516 15804
rect 7572 15802 7596 15804
rect 7652 15802 7658 15804
rect 7412 15750 7414 15802
rect 7594 15750 7596 15802
rect 7350 15748 7356 15750
rect 7412 15748 7436 15750
rect 7492 15748 7516 15750
rect 7572 15748 7596 15750
rect 7652 15748 7658 15750
rect 7350 15739 7658 15748
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14618 7236 14758
rect 7350 14716 7658 14725
rect 7350 14714 7356 14716
rect 7412 14714 7436 14716
rect 7492 14714 7516 14716
rect 7572 14714 7596 14716
rect 7652 14714 7658 14716
rect 7412 14662 7414 14714
rect 7594 14662 7596 14714
rect 7350 14660 7356 14662
rect 7412 14660 7436 14662
rect 7492 14660 7516 14662
rect 7572 14660 7596 14662
rect 7652 14660 7658 14662
rect 7350 14651 7658 14660
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7300 14006 7328 14486
rect 7852 14278 7880 15914
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7944 15570 7972 15846
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8010 15260 8318 15269
rect 8010 15258 8016 15260
rect 8072 15258 8096 15260
rect 8152 15258 8176 15260
rect 8232 15258 8256 15260
rect 8312 15258 8318 15260
rect 8072 15206 8074 15258
rect 8254 15206 8256 15258
rect 8010 15204 8016 15206
rect 8072 15204 8096 15206
rect 8152 15204 8176 15206
rect 8232 15204 8256 15206
rect 8312 15204 8318 15206
rect 8010 15195 8318 15204
rect 8404 15162 8432 15438
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8208 14816 8260 14822
rect 8864 14793 8892 14826
rect 8208 14758 8260 14764
rect 8850 14784 8906 14793
rect 8220 14482 8248 14758
rect 8850 14719 8906 14728
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7840 14272 7892 14278
rect 7760 14220 7840 14226
rect 7760 14214 7892 14220
rect 7760 14198 7880 14214
rect 7288 14000 7340 14006
rect 7208 13960 7288 13988
rect 7208 12986 7236 13960
rect 7288 13942 7340 13948
rect 7350 13628 7658 13637
rect 7350 13626 7356 13628
rect 7412 13626 7436 13628
rect 7492 13626 7516 13628
rect 7572 13626 7596 13628
rect 7652 13626 7658 13628
rect 7412 13574 7414 13626
rect 7594 13574 7596 13626
rect 7350 13572 7356 13574
rect 7412 13572 7436 13574
rect 7492 13572 7516 13574
rect 7572 13572 7596 13574
rect 7652 13572 7658 13574
rect 7350 13563 7658 13572
rect 7760 13274 7788 14198
rect 8010 14172 8318 14181
rect 8010 14170 8016 14172
rect 8072 14170 8096 14172
rect 8152 14170 8176 14172
rect 8232 14170 8256 14172
rect 8312 14170 8318 14172
rect 8072 14118 8074 14170
rect 8254 14118 8256 14170
rect 8010 14116 8016 14118
rect 8072 14116 8096 14118
rect 8152 14116 8176 14118
rect 8232 14116 8256 14118
rect 8312 14116 8318 14118
rect 8010 14107 8318 14116
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 13394 7880 13806
rect 8298 13424 8354 13433
rect 7840 13388 7892 13394
rect 8298 13359 8354 13368
rect 7840 13330 7892 13336
rect 7760 13246 7880 13274
rect 8312 13258 8340 13359
rect 7852 13190 7880 13246
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7116 12838 7236 12866
rect 7208 11778 7236 12838
rect 7350 12540 7658 12549
rect 7350 12538 7356 12540
rect 7412 12538 7436 12540
rect 7492 12538 7516 12540
rect 7572 12538 7596 12540
rect 7652 12538 7658 12540
rect 7412 12486 7414 12538
rect 7594 12486 7596 12538
rect 7350 12484 7356 12486
rect 7412 12484 7436 12486
rect 7492 12484 7516 12486
rect 7572 12484 7596 12486
rect 7652 12484 7658 12486
rect 7350 12475 7658 12484
rect 7852 12306 7880 13126
rect 8010 13084 8318 13093
rect 8010 13082 8016 13084
rect 8072 13082 8096 13084
rect 8152 13082 8176 13084
rect 8232 13082 8256 13084
rect 8312 13082 8318 13084
rect 8072 13030 8074 13082
rect 8254 13030 8256 13082
rect 8010 13028 8016 13030
rect 8072 13028 8096 13030
rect 8152 13028 8176 13030
rect 8232 13028 8256 13030
rect 8312 13028 8318 13030
rect 8010 13019 8318 13028
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8312 12434 8340 12582
rect 8312 12406 8432 12434
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7116 11750 7236 11778
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 9926 7052 10950
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 7993 7052 9522
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 7002 6960 7142
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7024 6934 7052 7686
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7116 6798 7144 11750
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7668 11642 7696 12038
rect 7760 11898 7788 12038
rect 7852 11898 7880 12038
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7944 11778 7972 12174
rect 8010 11996 8318 12005
rect 8010 11994 8016 11996
rect 8072 11994 8096 11996
rect 8152 11994 8176 11996
rect 8232 11994 8256 11996
rect 8312 11994 8318 11996
rect 8072 11942 8074 11994
rect 8254 11942 8256 11994
rect 8010 11940 8016 11942
rect 8072 11940 8096 11942
rect 8152 11940 8176 11942
rect 8232 11940 8256 11942
rect 8312 11940 8318 11942
rect 8010 11931 8318 11940
rect 7852 11750 7972 11778
rect 8404 11762 8432 12406
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8482 12064 8538 12073
rect 8482 11999 8538 12008
rect 8392 11756 8444 11762
rect 7208 11354 7236 11630
rect 7668 11614 7788 11642
rect 7350 11452 7658 11461
rect 7350 11450 7356 11452
rect 7412 11450 7436 11452
rect 7492 11450 7516 11452
rect 7572 11450 7596 11452
rect 7652 11450 7658 11452
rect 7412 11398 7414 11450
rect 7594 11398 7596 11450
rect 7350 11396 7356 11398
rect 7412 11396 7436 11398
rect 7492 11396 7516 11398
rect 7572 11396 7596 11398
rect 7652 11396 7658 11398
rect 7350 11387 7658 11396
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7760 10606 7788 11614
rect 7852 10690 7880 11750
rect 8392 11698 8444 11704
rect 8496 11694 8524 11999
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 10810 7972 11494
rect 8010 10908 8318 10917
rect 8010 10906 8016 10908
rect 8072 10906 8096 10908
rect 8152 10906 8176 10908
rect 8232 10906 8256 10908
rect 8312 10906 8318 10908
rect 8072 10854 8074 10906
rect 8254 10854 8256 10906
rect 8010 10852 8016 10854
rect 8072 10852 8096 10854
rect 8152 10852 8176 10854
rect 8232 10852 8256 10854
rect 8312 10852 8318 10854
rect 8010 10843 8318 10852
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7930 10704 7986 10713
rect 7852 10662 7930 10690
rect 7930 10639 7986 10648
rect 8588 10606 8616 12242
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10130 7236 10406
rect 7350 10364 7658 10373
rect 7350 10362 7356 10364
rect 7412 10362 7436 10364
rect 7492 10362 7516 10364
rect 7572 10362 7596 10364
rect 7652 10362 7658 10364
rect 7412 10310 7414 10362
rect 7594 10310 7596 10362
rect 7350 10308 7356 10310
rect 7412 10308 7436 10310
rect 7492 10308 7516 10310
rect 7572 10308 7596 10310
rect 7652 10308 7658 10310
rect 7350 10299 7658 10308
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7300 9674 7328 9930
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8010 9820 8318 9829
rect 8010 9818 8016 9820
rect 8072 9818 8096 9820
rect 8152 9818 8176 9820
rect 8232 9818 8256 9820
rect 8312 9818 8318 9820
rect 8072 9766 8074 9818
rect 8254 9766 8256 9818
rect 8010 9764 8016 9766
rect 8072 9764 8096 9766
rect 8152 9764 8176 9766
rect 8232 9764 8256 9766
rect 8312 9764 8318 9766
rect 8010 9755 8318 9764
rect 7208 9646 7328 9674
rect 7208 9058 7236 9646
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7350 9276 7658 9285
rect 7350 9274 7356 9276
rect 7412 9274 7436 9276
rect 7492 9274 7516 9276
rect 7572 9274 7596 9276
rect 7652 9274 7658 9276
rect 7412 9222 7414 9274
rect 7594 9222 7596 9274
rect 7350 9220 7356 9222
rect 7412 9220 7436 9222
rect 7492 9220 7516 9222
rect 7572 9220 7596 9222
rect 7652 9220 7658 9222
rect 7350 9211 7658 9220
rect 7760 9178 7788 9318
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7208 9030 7328 9058
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7208 8634 7236 8910
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7300 8566 7328 9030
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7288 8560 7340 8566
rect 7208 8508 7288 8514
rect 7208 8502 7340 8508
rect 7208 8486 7328 8502
rect 7208 7886 7236 8486
rect 7350 8188 7658 8197
rect 7350 8186 7356 8188
rect 7412 8186 7436 8188
rect 7492 8186 7516 8188
rect 7572 8186 7596 8188
rect 7652 8186 7658 8188
rect 7412 8134 7414 8186
rect 7594 8134 7596 8186
rect 7350 8132 7356 8134
rect 7412 8132 7436 8134
rect 7492 8132 7516 8134
rect 7572 8132 7596 8134
rect 7652 8132 7658 8134
rect 7350 8123 7658 8132
rect 7760 7886 7788 8774
rect 7852 7954 7880 9386
rect 7944 8090 7972 9386
rect 8128 9178 8156 9522
rect 8298 9344 8354 9353
rect 8298 9279 8354 9288
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8312 8974 8340 9279
rect 8404 9042 8432 9862
rect 8588 9518 8616 10542
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8010 8732 8318 8741
rect 8010 8730 8016 8732
rect 8072 8730 8096 8732
rect 8152 8730 8176 8732
rect 8232 8730 8256 8732
rect 8312 8730 8318 8732
rect 8072 8678 8074 8730
rect 8254 8678 8256 8730
rect 8010 8676 8016 8678
rect 8072 8676 8096 8678
rect 8152 8676 8176 8678
rect 8232 8676 8256 8678
rect 8312 8676 8318 8678
rect 8010 8667 8318 8676
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7748 7880 7800 7886
rect 7944 7834 7972 8026
rect 7748 7822 7800 7828
rect 7392 7478 7420 7822
rect 7852 7806 7972 7834
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7546 7788 7686
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7350 7100 7658 7109
rect 7350 7098 7356 7100
rect 7412 7098 7436 7100
rect 7492 7098 7516 7100
rect 7572 7098 7596 7100
rect 7652 7098 7658 7100
rect 7412 7046 7414 7098
rect 7594 7046 7596 7098
rect 7350 7044 7356 7046
rect 7412 7044 7436 7046
rect 7492 7044 7516 7046
rect 7572 7044 7596 7046
rect 7652 7044 7658 7046
rect 7350 7035 7658 7044
rect 7654 6896 7710 6905
rect 7852 6866 7880 7806
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7654 6831 7710 6840
rect 7840 6860 7892 6866
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2350 6012 2658 6021
rect 2350 6010 2356 6012
rect 2412 6010 2436 6012
rect 2492 6010 2516 6012
rect 2572 6010 2596 6012
rect 2652 6010 2658 6012
rect 2412 5958 2414 6010
rect 2594 5958 2596 6010
rect 2350 5956 2356 5958
rect 2412 5956 2436 5958
rect 2492 5956 2516 5958
rect 2572 5956 2596 5958
rect 2652 5956 2658 5958
rect 2350 5947 2658 5956
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2350 4924 2658 4933
rect 2350 4922 2356 4924
rect 2412 4922 2436 4924
rect 2492 4922 2516 4924
rect 2572 4922 2596 4924
rect 2652 4922 2658 4924
rect 2412 4870 2414 4922
rect 2594 4870 2596 4922
rect 2350 4868 2356 4870
rect 2412 4868 2436 4870
rect 2492 4868 2516 4870
rect 2572 4868 2596 4870
rect 2652 4868 2658 4870
rect 2350 4859 2658 4868
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2350 3836 2658 3845
rect 2350 3834 2356 3836
rect 2412 3834 2436 3836
rect 2492 3834 2516 3836
rect 2572 3834 2596 3836
rect 2652 3834 2658 3836
rect 2412 3782 2414 3834
rect 2594 3782 2596 3834
rect 2350 3780 2356 3782
rect 2412 3780 2436 3782
rect 2492 3780 2516 3782
rect 2572 3780 2596 3782
rect 2652 3780 2658 3782
rect 2350 3771 2658 3780
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 848 2848 900 2854
rect 848 2790 900 2796
rect 860 800 888 2790
rect 1872 2514 1900 2994
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 846 0 902 800
rect 2148 762 2176 2790
rect 2350 2748 2658 2757
rect 2350 2746 2356 2748
rect 2412 2746 2436 2748
rect 2492 2746 2516 2748
rect 2572 2746 2596 2748
rect 2652 2746 2658 2748
rect 2412 2694 2414 2746
rect 2594 2694 2596 2746
rect 2350 2692 2356 2694
rect 2412 2692 2436 2694
rect 2492 2692 2516 2694
rect 2572 2692 2596 2694
rect 2652 2692 2658 2694
rect 2350 2683 2658 2692
rect 5552 2446 5580 6598
rect 7116 6458 7144 6734
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7668 6390 7696 6831
rect 7840 6802 7892 6808
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6458 7880 6598
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7656 6384 7708 6390
rect 7708 6332 7788 6338
rect 7656 6326 7788 6332
rect 7668 6310 7788 6326
rect 7350 6012 7658 6021
rect 7350 6010 7356 6012
rect 7412 6010 7436 6012
rect 7492 6010 7516 6012
rect 7572 6010 7596 6012
rect 7652 6010 7658 6012
rect 7412 5958 7414 6010
rect 7594 5958 7596 6010
rect 7350 5956 7356 5958
rect 7412 5956 7436 5958
rect 7492 5956 7516 5958
rect 7572 5956 7596 5958
rect 7652 5956 7658 5958
rect 7350 5947 7658 5956
rect 7350 4924 7658 4933
rect 7350 4922 7356 4924
rect 7412 4922 7436 4924
rect 7492 4922 7516 4924
rect 7572 4922 7596 4924
rect 7652 4922 7658 4924
rect 7412 4870 7414 4922
rect 7594 4870 7596 4922
rect 7350 4868 7356 4870
rect 7412 4868 7436 4870
rect 7492 4868 7516 4870
rect 7572 4868 7596 4870
rect 7652 4868 7658 4870
rect 7350 4859 7658 4868
rect 7350 3836 7658 3845
rect 7350 3834 7356 3836
rect 7412 3834 7436 3836
rect 7492 3834 7516 3836
rect 7572 3834 7596 3836
rect 7652 3834 7658 3836
rect 7412 3782 7414 3834
rect 7594 3782 7596 3834
rect 7350 3780 7356 3782
rect 7412 3780 7436 3782
rect 7492 3780 7516 3782
rect 7572 3780 7596 3782
rect 7652 3780 7658 3782
rect 7350 3771 7658 3780
rect 7350 2748 7658 2757
rect 7350 2746 7356 2748
rect 7412 2746 7436 2748
rect 7492 2746 7516 2748
rect 7572 2746 7596 2748
rect 7652 2746 7658 2748
rect 7412 2694 7414 2746
rect 7594 2694 7596 2746
rect 7350 2692 7356 2694
rect 7412 2692 7436 2694
rect 7492 2692 7516 2694
rect 7572 2692 7596 2694
rect 7652 2692 7658 2694
rect 6642 2680 6698 2689
rect 7350 2683 7658 2692
rect 7760 2650 7788 6310
rect 7944 2650 7972 7686
rect 8010 7644 8318 7653
rect 8010 7642 8016 7644
rect 8072 7642 8096 7644
rect 8152 7642 8176 7644
rect 8232 7642 8256 7644
rect 8312 7642 8318 7644
rect 8072 7590 8074 7642
rect 8254 7590 8256 7642
rect 8010 7588 8016 7590
rect 8072 7588 8096 7590
rect 8152 7588 8176 7590
rect 8232 7588 8256 7590
rect 8312 7588 8318 7590
rect 8010 7579 8318 7588
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8010 6556 8318 6565
rect 8010 6554 8016 6556
rect 8072 6554 8096 6556
rect 8152 6554 8176 6556
rect 8232 6554 8256 6556
rect 8312 6554 8318 6556
rect 8072 6502 8074 6554
rect 8254 6502 8256 6554
rect 8010 6500 8016 6502
rect 8072 6500 8096 6502
rect 8152 6500 8176 6502
rect 8232 6500 8256 6502
rect 8312 6500 8318 6502
rect 8010 6491 8318 6500
rect 8404 6322 8432 7142
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8850 6624 8906 6633
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8496 5914 8524 6598
rect 8850 6559 8906 6568
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8864 5710 8892 6559
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8010 5468 8318 5477
rect 8010 5466 8016 5468
rect 8072 5466 8096 5468
rect 8152 5466 8176 5468
rect 8232 5466 8256 5468
rect 8312 5466 8318 5468
rect 8072 5414 8074 5466
rect 8254 5414 8256 5466
rect 8010 5412 8016 5414
rect 8072 5412 8096 5414
rect 8152 5412 8176 5414
rect 8232 5412 8256 5414
rect 8312 5412 8318 5414
rect 8010 5403 8318 5412
rect 8010 4380 8318 4389
rect 8010 4378 8016 4380
rect 8072 4378 8096 4380
rect 8152 4378 8176 4380
rect 8232 4378 8256 4380
rect 8312 4378 8318 4380
rect 8072 4326 8074 4378
rect 8254 4326 8256 4378
rect 8010 4324 8016 4326
rect 8072 4324 8096 4326
rect 8152 4324 8176 4326
rect 8232 4324 8256 4326
rect 8312 4324 8318 4326
rect 8010 4315 8318 4324
rect 8010 3292 8318 3301
rect 8010 3290 8016 3292
rect 8072 3290 8096 3292
rect 8152 3290 8176 3292
rect 8232 3290 8256 3292
rect 8312 3290 8318 3292
rect 8072 3238 8074 3290
rect 8254 3238 8256 3290
rect 8010 3236 8016 3238
rect 8072 3236 8096 3238
rect 8152 3236 8176 3238
rect 8232 3236 8256 3238
rect 8312 3236 8318 3238
rect 8010 3227 8318 3236
rect 6642 2615 6698 2624
rect 7748 2644 7800 2650
rect 6656 2514 6684 2615
rect 7748 2586 7800 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2424 870 2544 898
rect 2424 762 2452 870
rect 2516 800 2544 870
rect 4172 800 4200 2246
rect 5828 800 5856 2382
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 7668 1170 7696 2314
rect 8010 2204 8318 2213
rect 8010 2202 8016 2204
rect 8072 2202 8096 2204
rect 8152 2202 8176 2204
rect 8232 2202 8256 2204
rect 8312 2202 8318 2204
rect 8072 2150 8074 2202
rect 8254 2150 8256 2202
rect 8010 2148 8016 2150
rect 8072 2148 8096 2150
rect 8152 2148 8176 2150
rect 8232 2148 8256 2150
rect 8312 2148 8318 2150
rect 8010 2139 8318 2148
rect 7484 1142 7696 1170
rect 7484 800 7512 1142
rect 9140 800 9168 2314
rect 2148 734 2452 762
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7470 0 7526 800
rect 9126 0 9182 800
<< via2 >>
rect 2356 77818 2412 77820
rect 2436 77818 2492 77820
rect 2516 77818 2572 77820
rect 2596 77818 2652 77820
rect 2356 77766 2402 77818
rect 2402 77766 2412 77818
rect 2436 77766 2466 77818
rect 2466 77766 2478 77818
rect 2478 77766 2492 77818
rect 2516 77766 2530 77818
rect 2530 77766 2542 77818
rect 2542 77766 2572 77818
rect 2596 77766 2606 77818
rect 2606 77766 2652 77818
rect 2356 77764 2412 77766
rect 2436 77764 2492 77766
rect 2516 77764 2572 77766
rect 2596 77764 2652 77766
rect 3016 77274 3072 77276
rect 3096 77274 3152 77276
rect 3176 77274 3232 77276
rect 3256 77274 3312 77276
rect 3016 77222 3062 77274
rect 3062 77222 3072 77274
rect 3096 77222 3126 77274
rect 3126 77222 3138 77274
rect 3138 77222 3152 77274
rect 3176 77222 3190 77274
rect 3190 77222 3202 77274
rect 3202 77222 3232 77274
rect 3256 77222 3266 77274
rect 3266 77222 3312 77274
rect 3016 77220 3072 77222
rect 3096 77220 3152 77222
rect 3176 77220 3232 77222
rect 3256 77220 3312 77222
rect 2356 76730 2412 76732
rect 2436 76730 2492 76732
rect 2516 76730 2572 76732
rect 2596 76730 2652 76732
rect 2356 76678 2402 76730
rect 2402 76678 2412 76730
rect 2436 76678 2466 76730
rect 2466 76678 2478 76730
rect 2478 76678 2492 76730
rect 2516 76678 2530 76730
rect 2530 76678 2542 76730
rect 2542 76678 2572 76730
rect 2596 76678 2606 76730
rect 2606 76678 2652 76730
rect 2356 76676 2412 76678
rect 2436 76676 2492 76678
rect 2516 76676 2572 76678
rect 2596 76676 2652 76678
rect 3016 76186 3072 76188
rect 3096 76186 3152 76188
rect 3176 76186 3232 76188
rect 3256 76186 3312 76188
rect 3016 76134 3062 76186
rect 3062 76134 3072 76186
rect 3096 76134 3126 76186
rect 3126 76134 3138 76186
rect 3138 76134 3152 76186
rect 3176 76134 3190 76186
rect 3190 76134 3202 76186
rect 3202 76134 3232 76186
rect 3256 76134 3266 76186
rect 3266 76134 3312 76186
rect 3016 76132 3072 76134
rect 3096 76132 3152 76134
rect 3176 76132 3232 76134
rect 3256 76132 3312 76134
rect 2356 75642 2412 75644
rect 2436 75642 2492 75644
rect 2516 75642 2572 75644
rect 2596 75642 2652 75644
rect 2356 75590 2402 75642
rect 2402 75590 2412 75642
rect 2436 75590 2466 75642
rect 2466 75590 2478 75642
rect 2478 75590 2492 75642
rect 2516 75590 2530 75642
rect 2530 75590 2542 75642
rect 2542 75590 2572 75642
rect 2596 75590 2606 75642
rect 2606 75590 2652 75642
rect 2356 75588 2412 75590
rect 2436 75588 2492 75590
rect 2516 75588 2572 75590
rect 2596 75588 2652 75590
rect 3016 75098 3072 75100
rect 3096 75098 3152 75100
rect 3176 75098 3232 75100
rect 3256 75098 3312 75100
rect 3016 75046 3062 75098
rect 3062 75046 3072 75098
rect 3096 75046 3126 75098
rect 3126 75046 3138 75098
rect 3138 75046 3152 75098
rect 3176 75046 3190 75098
rect 3190 75046 3202 75098
rect 3202 75046 3232 75098
rect 3256 75046 3266 75098
rect 3266 75046 3312 75098
rect 3016 75044 3072 75046
rect 3096 75044 3152 75046
rect 3176 75044 3232 75046
rect 3256 75044 3312 75046
rect 2356 74554 2412 74556
rect 2436 74554 2492 74556
rect 2516 74554 2572 74556
rect 2596 74554 2652 74556
rect 2356 74502 2402 74554
rect 2402 74502 2412 74554
rect 2436 74502 2466 74554
rect 2466 74502 2478 74554
rect 2478 74502 2492 74554
rect 2516 74502 2530 74554
rect 2530 74502 2542 74554
rect 2542 74502 2572 74554
rect 2596 74502 2606 74554
rect 2606 74502 2652 74554
rect 2356 74500 2412 74502
rect 2436 74500 2492 74502
rect 2516 74500 2572 74502
rect 2596 74500 2652 74502
rect 3016 74010 3072 74012
rect 3096 74010 3152 74012
rect 3176 74010 3232 74012
rect 3256 74010 3312 74012
rect 3016 73958 3062 74010
rect 3062 73958 3072 74010
rect 3096 73958 3126 74010
rect 3126 73958 3138 74010
rect 3138 73958 3152 74010
rect 3176 73958 3190 74010
rect 3190 73958 3202 74010
rect 3202 73958 3232 74010
rect 3256 73958 3266 74010
rect 3266 73958 3312 74010
rect 3016 73956 3072 73958
rect 3096 73956 3152 73958
rect 3176 73956 3232 73958
rect 3256 73956 3312 73958
rect 2356 73466 2412 73468
rect 2436 73466 2492 73468
rect 2516 73466 2572 73468
rect 2596 73466 2652 73468
rect 2356 73414 2402 73466
rect 2402 73414 2412 73466
rect 2436 73414 2466 73466
rect 2466 73414 2478 73466
rect 2478 73414 2492 73466
rect 2516 73414 2530 73466
rect 2530 73414 2542 73466
rect 2542 73414 2572 73466
rect 2596 73414 2606 73466
rect 2606 73414 2652 73466
rect 2356 73412 2412 73414
rect 2436 73412 2492 73414
rect 2516 73412 2572 73414
rect 2596 73412 2652 73414
rect 3016 72922 3072 72924
rect 3096 72922 3152 72924
rect 3176 72922 3232 72924
rect 3256 72922 3312 72924
rect 3016 72870 3062 72922
rect 3062 72870 3072 72922
rect 3096 72870 3126 72922
rect 3126 72870 3138 72922
rect 3138 72870 3152 72922
rect 3176 72870 3190 72922
rect 3190 72870 3202 72922
rect 3202 72870 3232 72922
rect 3256 72870 3266 72922
rect 3266 72870 3312 72922
rect 3016 72868 3072 72870
rect 3096 72868 3152 72870
rect 3176 72868 3232 72870
rect 3256 72868 3312 72870
rect 2356 72378 2412 72380
rect 2436 72378 2492 72380
rect 2516 72378 2572 72380
rect 2596 72378 2652 72380
rect 2356 72326 2402 72378
rect 2402 72326 2412 72378
rect 2436 72326 2466 72378
rect 2466 72326 2478 72378
rect 2478 72326 2492 72378
rect 2516 72326 2530 72378
rect 2530 72326 2542 72378
rect 2542 72326 2572 72378
rect 2596 72326 2606 72378
rect 2606 72326 2652 72378
rect 2356 72324 2412 72326
rect 2436 72324 2492 72326
rect 2516 72324 2572 72326
rect 2596 72324 2652 72326
rect 3016 71834 3072 71836
rect 3096 71834 3152 71836
rect 3176 71834 3232 71836
rect 3256 71834 3312 71836
rect 3016 71782 3062 71834
rect 3062 71782 3072 71834
rect 3096 71782 3126 71834
rect 3126 71782 3138 71834
rect 3138 71782 3152 71834
rect 3176 71782 3190 71834
rect 3190 71782 3202 71834
rect 3202 71782 3232 71834
rect 3256 71782 3266 71834
rect 3266 71782 3312 71834
rect 3016 71780 3072 71782
rect 3096 71780 3152 71782
rect 3176 71780 3232 71782
rect 3256 71780 3312 71782
rect 2356 71290 2412 71292
rect 2436 71290 2492 71292
rect 2516 71290 2572 71292
rect 2596 71290 2652 71292
rect 2356 71238 2402 71290
rect 2402 71238 2412 71290
rect 2436 71238 2466 71290
rect 2466 71238 2478 71290
rect 2478 71238 2492 71290
rect 2516 71238 2530 71290
rect 2530 71238 2542 71290
rect 2542 71238 2572 71290
rect 2596 71238 2606 71290
rect 2606 71238 2652 71290
rect 2356 71236 2412 71238
rect 2436 71236 2492 71238
rect 2516 71236 2572 71238
rect 2596 71236 2652 71238
rect 3016 70746 3072 70748
rect 3096 70746 3152 70748
rect 3176 70746 3232 70748
rect 3256 70746 3312 70748
rect 3016 70694 3062 70746
rect 3062 70694 3072 70746
rect 3096 70694 3126 70746
rect 3126 70694 3138 70746
rect 3138 70694 3152 70746
rect 3176 70694 3190 70746
rect 3190 70694 3202 70746
rect 3202 70694 3232 70746
rect 3256 70694 3266 70746
rect 3266 70694 3312 70746
rect 3016 70692 3072 70694
rect 3096 70692 3152 70694
rect 3176 70692 3232 70694
rect 3256 70692 3312 70694
rect 2356 70202 2412 70204
rect 2436 70202 2492 70204
rect 2516 70202 2572 70204
rect 2596 70202 2652 70204
rect 2356 70150 2402 70202
rect 2402 70150 2412 70202
rect 2436 70150 2466 70202
rect 2466 70150 2478 70202
rect 2478 70150 2492 70202
rect 2516 70150 2530 70202
rect 2530 70150 2542 70202
rect 2542 70150 2572 70202
rect 2596 70150 2606 70202
rect 2606 70150 2652 70202
rect 2356 70148 2412 70150
rect 2436 70148 2492 70150
rect 2516 70148 2572 70150
rect 2596 70148 2652 70150
rect 3016 69658 3072 69660
rect 3096 69658 3152 69660
rect 3176 69658 3232 69660
rect 3256 69658 3312 69660
rect 3016 69606 3062 69658
rect 3062 69606 3072 69658
rect 3096 69606 3126 69658
rect 3126 69606 3138 69658
rect 3138 69606 3152 69658
rect 3176 69606 3190 69658
rect 3190 69606 3202 69658
rect 3202 69606 3232 69658
rect 3256 69606 3266 69658
rect 3266 69606 3312 69658
rect 3016 69604 3072 69606
rect 3096 69604 3152 69606
rect 3176 69604 3232 69606
rect 3256 69604 3312 69606
rect 2356 69114 2412 69116
rect 2436 69114 2492 69116
rect 2516 69114 2572 69116
rect 2596 69114 2652 69116
rect 2356 69062 2402 69114
rect 2402 69062 2412 69114
rect 2436 69062 2466 69114
rect 2466 69062 2478 69114
rect 2478 69062 2492 69114
rect 2516 69062 2530 69114
rect 2530 69062 2542 69114
rect 2542 69062 2572 69114
rect 2596 69062 2606 69114
rect 2606 69062 2652 69114
rect 2356 69060 2412 69062
rect 2436 69060 2492 69062
rect 2516 69060 2572 69062
rect 2596 69060 2652 69062
rect 3016 68570 3072 68572
rect 3096 68570 3152 68572
rect 3176 68570 3232 68572
rect 3256 68570 3312 68572
rect 3016 68518 3062 68570
rect 3062 68518 3072 68570
rect 3096 68518 3126 68570
rect 3126 68518 3138 68570
rect 3138 68518 3152 68570
rect 3176 68518 3190 68570
rect 3190 68518 3202 68570
rect 3202 68518 3232 68570
rect 3256 68518 3266 68570
rect 3266 68518 3312 68570
rect 3016 68516 3072 68518
rect 3096 68516 3152 68518
rect 3176 68516 3232 68518
rect 3256 68516 3312 68518
rect 2356 68026 2412 68028
rect 2436 68026 2492 68028
rect 2516 68026 2572 68028
rect 2596 68026 2652 68028
rect 2356 67974 2402 68026
rect 2402 67974 2412 68026
rect 2436 67974 2466 68026
rect 2466 67974 2478 68026
rect 2478 67974 2492 68026
rect 2516 67974 2530 68026
rect 2530 67974 2542 68026
rect 2542 67974 2572 68026
rect 2596 67974 2606 68026
rect 2606 67974 2652 68026
rect 2356 67972 2412 67974
rect 2436 67972 2492 67974
rect 2516 67972 2572 67974
rect 2596 67972 2652 67974
rect 3016 67482 3072 67484
rect 3096 67482 3152 67484
rect 3176 67482 3232 67484
rect 3256 67482 3312 67484
rect 3016 67430 3062 67482
rect 3062 67430 3072 67482
rect 3096 67430 3126 67482
rect 3126 67430 3138 67482
rect 3138 67430 3152 67482
rect 3176 67430 3190 67482
rect 3190 67430 3202 67482
rect 3202 67430 3232 67482
rect 3256 67430 3266 67482
rect 3266 67430 3312 67482
rect 3016 67428 3072 67430
rect 3096 67428 3152 67430
rect 3176 67428 3232 67430
rect 3256 67428 3312 67430
rect 2356 66938 2412 66940
rect 2436 66938 2492 66940
rect 2516 66938 2572 66940
rect 2596 66938 2652 66940
rect 2356 66886 2402 66938
rect 2402 66886 2412 66938
rect 2436 66886 2466 66938
rect 2466 66886 2478 66938
rect 2478 66886 2492 66938
rect 2516 66886 2530 66938
rect 2530 66886 2542 66938
rect 2542 66886 2572 66938
rect 2596 66886 2606 66938
rect 2606 66886 2652 66938
rect 2356 66884 2412 66886
rect 2436 66884 2492 66886
rect 2516 66884 2572 66886
rect 2596 66884 2652 66886
rect 3016 66394 3072 66396
rect 3096 66394 3152 66396
rect 3176 66394 3232 66396
rect 3256 66394 3312 66396
rect 3016 66342 3062 66394
rect 3062 66342 3072 66394
rect 3096 66342 3126 66394
rect 3126 66342 3138 66394
rect 3138 66342 3152 66394
rect 3176 66342 3190 66394
rect 3190 66342 3202 66394
rect 3202 66342 3232 66394
rect 3256 66342 3266 66394
rect 3266 66342 3312 66394
rect 3016 66340 3072 66342
rect 3096 66340 3152 66342
rect 3176 66340 3232 66342
rect 3256 66340 3312 66342
rect 2356 65850 2412 65852
rect 2436 65850 2492 65852
rect 2516 65850 2572 65852
rect 2596 65850 2652 65852
rect 2356 65798 2402 65850
rect 2402 65798 2412 65850
rect 2436 65798 2466 65850
rect 2466 65798 2478 65850
rect 2478 65798 2492 65850
rect 2516 65798 2530 65850
rect 2530 65798 2542 65850
rect 2542 65798 2572 65850
rect 2596 65798 2606 65850
rect 2606 65798 2652 65850
rect 2356 65796 2412 65798
rect 2436 65796 2492 65798
rect 2516 65796 2572 65798
rect 2596 65796 2652 65798
rect 3016 65306 3072 65308
rect 3096 65306 3152 65308
rect 3176 65306 3232 65308
rect 3256 65306 3312 65308
rect 3016 65254 3062 65306
rect 3062 65254 3072 65306
rect 3096 65254 3126 65306
rect 3126 65254 3138 65306
rect 3138 65254 3152 65306
rect 3176 65254 3190 65306
rect 3190 65254 3202 65306
rect 3202 65254 3232 65306
rect 3256 65254 3266 65306
rect 3266 65254 3312 65306
rect 3016 65252 3072 65254
rect 3096 65252 3152 65254
rect 3176 65252 3232 65254
rect 3256 65252 3312 65254
rect 2356 64762 2412 64764
rect 2436 64762 2492 64764
rect 2516 64762 2572 64764
rect 2596 64762 2652 64764
rect 2356 64710 2402 64762
rect 2402 64710 2412 64762
rect 2436 64710 2466 64762
rect 2466 64710 2478 64762
rect 2478 64710 2492 64762
rect 2516 64710 2530 64762
rect 2530 64710 2542 64762
rect 2542 64710 2572 64762
rect 2596 64710 2606 64762
rect 2606 64710 2652 64762
rect 2356 64708 2412 64710
rect 2436 64708 2492 64710
rect 2516 64708 2572 64710
rect 2596 64708 2652 64710
rect 3016 64218 3072 64220
rect 3096 64218 3152 64220
rect 3176 64218 3232 64220
rect 3256 64218 3312 64220
rect 3016 64166 3062 64218
rect 3062 64166 3072 64218
rect 3096 64166 3126 64218
rect 3126 64166 3138 64218
rect 3138 64166 3152 64218
rect 3176 64166 3190 64218
rect 3190 64166 3202 64218
rect 3202 64166 3232 64218
rect 3256 64166 3266 64218
rect 3266 64166 3312 64218
rect 3016 64164 3072 64166
rect 3096 64164 3152 64166
rect 3176 64164 3232 64166
rect 3256 64164 3312 64166
rect 2356 63674 2412 63676
rect 2436 63674 2492 63676
rect 2516 63674 2572 63676
rect 2596 63674 2652 63676
rect 2356 63622 2402 63674
rect 2402 63622 2412 63674
rect 2436 63622 2466 63674
rect 2466 63622 2478 63674
rect 2478 63622 2492 63674
rect 2516 63622 2530 63674
rect 2530 63622 2542 63674
rect 2542 63622 2572 63674
rect 2596 63622 2606 63674
rect 2606 63622 2652 63674
rect 2356 63620 2412 63622
rect 2436 63620 2492 63622
rect 2516 63620 2572 63622
rect 2596 63620 2652 63622
rect 3016 63130 3072 63132
rect 3096 63130 3152 63132
rect 3176 63130 3232 63132
rect 3256 63130 3312 63132
rect 3016 63078 3062 63130
rect 3062 63078 3072 63130
rect 3096 63078 3126 63130
rect 3126 63078 3138 63130
rect 3138 63078 3152 63130
rect 3176 63078 3190 63130
rect 3190 63078 3202 63130
rect 3202 63078 3232 63130
rect 3256 63078 3266 63130
rect 3266 63078 3312 63130
rect 3016 63076 3072 63078
rect 3096 63076 3152 63078
rect 3176 63076 3232 63078
rect 3256 63076 3312 63078
rect 2356 62586 2412 62588
rect 2436 62586 2492 62588
rect 2516 62586 2572 62588
rect 2596 62586 2652 62588
rect 2356 62534 2402 62586
rect 2402 62534 2412 62586
rect 2436 62534 2466 62586
rect 2466 62534 2478 62586
rect 2478 62534 2492 62586
rect 2516 62534 2530 62586
rect 2530 62534 2542 62586
rect 2542 62534 2572 62586
rect 2596 62534 2606 62586
rect 2606 62534 2652 62586
rect 2356 62532 2412 62534
rect 2436 62532 2492 62534
rect 2516 62532 2572 62534
rect 2596 62532 2652 62534
rect 3016 62042 3072 62044
rect 3096 62042 3152 62044
rect 3176 62042 3232 62044
rect 3256 62042 3312 62044
rect 3016 61990 3062 62042
rect 3062 61990 3072 62042
rect 3096 61990 3126 62042
rect 3126 61990 3138 62042
rect 3138 61990 3152 62042
rect 3176 61990 3190 62042
rect 3190 61990 3202 62042
rect 3202 61990 3232 62042
rect 3256 61990 3266 62042
rect 3266 61990 3312 62042
rect 3016 61988 3072 61990
rect 3096 61988 3152 61990
rect 3176 61988 3232 61990
rect 3256 61988 3312 61990
rect 2356 61498 2412 61500
rect 2436 61498 2492 61500
rect 2516 61498 2572 61500
rect 2596 61498 2652 61500
rect 2356 61446 2402 61498
rect 2402 61446 2412 61498
rect 2436 61446 2466 61498
rect 2466 61446 2478 61498
rect 2478 61446 2492 61498
rect 2516 61446 2530 61498
rect 2530 61446 2542 61498
rect 2542 61446 2572 61498
rect 2596 61446 2606 61498
rect 2606 61446 2652 61498
rect 2356 61444 2412 61446
rect 2436 61444 2492 61446
rect 2516 61444 2572 61446
rect 2596 61444 2652 61446
rect 3016 60954 3072 60956
rect 3096 60954 3152 60956
rect 3176 60954 3232 60956
rect 3256 60954 3312 60956
rect 3016 60902 3062 60954
rect 3062 60902 3072 60954
rect 3096 60902 3126 60954
rect 3126 60902 3138 60954
rect 3138 60902 3152 60954
rect 3176 60902 3190 60954
rect 3190 60902 3202 60954
rect 3202 60902 3232 60954
rect 3256 60902 3266 60954
rect 3266 60902 3312 60954
rect 3016 60900 3072 60902
rect 3096 60900 3152 60902
rect 3176 60900 3232 60902
rect 3256 60900 3312 60902
rect 2356 60410 2412 60412
rect 2436 60410 2492 60412
rect 2516 60410 2572 60412
rect 2596 60410 2652 60412
rect 2356 60358 2402 60410
rect 2402 60358 2412 60410
rect 2436 60358 2466 60410
rect 2466 60358 2478 60410
rect 2478 60358 2492 60410
rect 2516 60358 2530 60410
rect 2530 60358 2542 60410
rect 2542 60358 2572 60410
rect 2596 60358 2606 60410
rect 2606 60358 2652 60410
rect 2356 60356 2412 60358
rect 2436 60356 2492 60358
rect 2516 60356 2572 60358
rect 2596 60356 2652 60358
rect 3016 59866 3072 59868
rect 3096 59866 3152 59868
rect 3176 59866 3232 59868
rect 3256 59866 3312 59868
rect 3016 59814 3062 59866
rect 3062 59814 3072 59866
rect 3096 59814 3126 59866
rect 3126 59814 3138 59866
rect 3138 59814 3152 59866
rect 3176 59814 3190 59866
rect 3190 59814 3202 59866
rect 3202 59814 3232 59866
rect 3256 59814 3266 59866
rect 3266 59814 3312 59866
rect 3016 59812 3072 59814
rect 3096 59812 3152 59814
rect 3176 59812 3232 59814
rect 3256 59812 3312 59814
rect 2356 59322 2412 59324
rect 2436 59322 2492 59324
rect 2516 59322 2572 59324
rect 2596 59322 2652 59324
rect 2356 59270 2402 59322
rect 2402 59270 2412 59322
rect 2436 59270 2466 59322
rect 2466 59270 2478 59322
rect 2478 59270 2492 59322
rect 2516 59270 2530 59322
rect 2530 59270 2542 59322
rect 2542 59270 2572 59322
rect 2596 59270 2606 59322
rect 2606 59270 2652 59322
rect 2356 59268 2412 59270
rect 2436 59268 2492 59270
rect 2516 59268 2572 59270
rect 2596 59268 2652 59270
rect 3016 58778 3072 58780
rect 3096 58778 3152 58780
rect 3176 58778 3232 58780
rect 3256 58778 3312 58780
rect 3016 58726 3062 58778
rect 3062 58726 3072 58778
rect 3096 58726 3126 58778
rect 3126 58726 3138 58778
rect 3138 58726 3152 58778
rect 3176 58726 3190 58778
rect 3190 58726 3202 58778
rect 3202 58726 3232 58778
rect 3256 58726 3266 58778
rect 3266 58726 3312 58778
rect 3016 58724 3072 58726
rect 3096 58724 3152 58726
rect 3176 58724 3232 58726
rect 3256 58724 3312 58726
rect 2356 58234 2412 58236
rect 2436 58234 2492 58236
rect 2516 58234 2572 58236
rect 2596 58234 2652 58236
rect 2356 58182 2402 58234
rect 2402 58182 2412 58234
rect 2436 58182 2466 58234
rect 2466 58182 2478 58234
rect 2478 58182 2492 58234
rect 2516 58182 2530 58234
rect 2530 58182 2542 58234
rect 2542 58182 2572 58234
rect 2596 58182 2606 58234
rect 2606 58182 2652 58234
rect 2356 58180 2412 58182
rect 2436 58180 2492 58182
rect 2516 58180 2572 58182
rect 2596 58180 2652 58182
rect 3016 57690 3072 57692
rect 3096 57690 3152 57692
rect 3176 57690 3232 57692
rect 3256 57690 3312 57692
rect 3016 57638 3062 57690
rect 3062 57638 3072 57690
rect 3096 57638 3126 57690
rect 3126 57638 3138 57690
rect 3138 57638 3152 57690
rect 3176 57638 3190 57690
rect 3190 57638 3202 57690
rect 3202 57638 3232 57690
rect 3256 57638 3266 57690
rect 3266 57638 3312 57690
rect 3016 57636 3072 57638
rect 3096 57636 3152 57638
rect 3176 57636 3232 57638
rect 3256 57636 3312 57638
rect 2356 57146 2412 57148
rect 2436 57146 2492 57148
rect 2516 57146 2572 57148
rect 2596 57146 2652 57148
rect 2356 57094 2402 57146
rect 2402 57094 2412 57146
rect 2436 57094 2466 57146
rect 2466 57094 2478 57146
rect 2478 57094 2492 57146
rect 2516 57094 2530 57146
rect 2530 57094 2542 57146
rect 2542 57094 2572 57146
rect 2596 57094 2606 57146
rect 2606 57094 2652 57146
rect 2356 57092 2412 57094
rect 2436 57092 2492 57094
rect 2516 57092 2572 57094
rect 2596 57092 2652 57094
rect 3016 56602 3072 56604
rect 3096 56602 3152 56604
rect 3176 56602 3232 56604
rect 3256 56602 3312 56604
rect 3016 56550 3062 56602
rect 3062 56550 3072 56602
rect 3096 56550 3126 56602
rect 3126 56550 3138 56602
rect 3138 56550 3152 56602
rect 3176 56550 3190 56602
rect 3190 56550 3202 56602
rect 3202 56550 3232 56602
rect 3256 56550 3266 56602
rect 3266 56550 3312 56602
rect 3016 56548 3072 56550
rect 3096 56548 3152 56550
rect 3176 56548 3232 56550
rect 3256 56548 3312 56550
rect 2356 56058 2412 56060
rect 2436 56058 2492 56060
rect 2516 56058 2572 56060
rect 2596 56058 2652 56060
rect 2356 56006 2402 56058
rect 2402 56006 2412 56058
rect 2436 56006 2466 56058
rect 2466 56006 2478 56058
rect 2478 56006 2492 56058
rect 2516 56006 2530 56058
rect 2530 56006 2542 56058
rect 2542 56006 2572 56058
rect 2596 56006 2606 56058
rect 2606 56006 2652 56058
rect 2356 56004 2412 56006
rect 2436 56004 2492 56006
rect 2516 56004 2572 56006
rect 2596 56004 2652 56006
rect 3016 55514 3072 55516
rect 3096 55514 3152 55516
rect 3176 55514 3232 55516
rect 3256 55514 3312 55516
rect 3016 55462 3062 55514
rect 3062 55462 3072 55514
rect 3096 55462 3126 55514
rect 3126 55462 3138 55514
rect 3138 55462 3152 55514
rect 3176 55462 3190 55514
rect 3190 55462 3202 55514
rect 3202 55462 3232 55514
rect 3256 55462 3266 55514
rect 3266 55462 3312 55514
rect 3016 55460 3072 55462
rect 3096 55460 3152 55462
rect 3176 55460 3232 55462
rect 3256 55460 3312 55462
rect 2356 54970 2412 54972
rect 2436 54970 2492 54972
rect 2516 54970 2572 54972
rect 2596 54970 2652 54972
rect 2356 54918 2402 54970
rect 2402 54918 2412 54970
rect 2436 54918 2466 54970
rect 2466 54918 2478 54970
rect 2478 54918 2492 54970
rect 2516 54918 2530 54970
rect 2530 54918 2542 54970
rect 2542 54918 2572 54970
rect 2596 54918 2606 54970
rect 2606 54918 2652 54970
rect 2356 54916 2412 54918
rect 2436 54916 2492 54918
rect 2516 54916 2572 54918
rect 2596 54916 2652 54918
rect 3016 54426 3072 54428
rect 3096 54426 3152 54428
rect 3176 54426 3232 54428
rect 3256 54426 3312 54428
rect 3016 54374 3062 54426
rect 3062 54374 3072 54426
rect 3096 54374 3126 54426
rect 3126 54374 3138 54426
rect 3138 54374 3152 54426
rect 3176 54374 3190 54426
rect 3190 54374 3202 54426
rect 3202 54374 3232 54426
rect 3256 54374 3266 54426
rect 3266 54374 3312 54426
rect 3016 54372 3072 54374
rect 3096 54372 3152 54374
rect 3176 54372 3232 54374
rect 3256 54372 3312 54374
rect 2356 53882 2412 53884
rect 2436 53882 2492 53884
rect 2516 53882 2572 53884
rect 2596 53882 2652 53884
rect 2356 53830 2402 53882
rect 2402 53830 2412 53882
rect 2436 53830 2466 53882
rect 2466 53830 2478 53882
rect 2478 53830 2492 53882
rect 2516 53830 2530 53882
rect 2530 53830 2542 53882
rect 2542 53830 2572 53882
rect 2596 53830 2606 53882
rect 2606 53830 2652 53882
rect 2356 53828 2412 53830
rect 2436 53828 2492 53830
rect 2516 53828 2572 53830
rect 2596 53828 2652 53830
rect 3016 53338 3072 53340
rect 3096 53338 3152 53340
rect 3176 53338 3232 53340
rect 3256 53338 3312 53340
rect 3016 53286 3062 53338
rect 3062 53286 3072 53338
rect 3096 53286 3126 53338
rect 3126 53286 3138 53338
rect 3138 53286 3152 53338
rect 3176 53286 3190 53338
rect 3190 53286 3202 53338
rect 3202 53286 3232 53338
rect 3256 53286 3266 53338
rect 3266 53286 3312 53338
rect 3016 53284 3072 53286
rect 3096 53284 3152 53286
rect 3176 53284 3232 53286
rect 3256 53284 3312 53286
rect 2356 52794 2412 52796
rect 2436 52794 2492 52796
rect 2516 52794 2572 52796
rect 2596 52794 2652 52796
rect 2356 52742 2402 52794
rect 2402 52742 2412 52794
rect 2436 52742 2466 52794
rect 2466 52742 2478 52794
rect 2478 52742 2492 52794
rect 2516 52742 2530 52794
rect 2530 52742 2542 52794
rect 2542 52742 2572 52794
rect 2596 52742 2606 52794
rect 2606 52742 2652 52794
rect 2356 52740 2412 52742
rect 2436 52740 2492 52742
rect 2516 52740 2572 52742
rect 2596 52740 2652 52742
rect 3016 52250 3072 52252
rect 3096 52250 3152 52252
rect 3176 52250 3232 52252
rect 3256 52250 3312 52252
rect 3016 52198 3062 52250
rect 3062 52198 3072 52250
rect 3096 52198 3126 52250
rect 3126 52198 3138 52250
rect 3138 52198 3152 52250
rect 3176 52198 3190 52250
rect 3190 52198 3202 52250
rect 3202 52198 3232 52250
rect 3256 52198 3266 52250
rect 3266 52198 3312 52250
rect 3016 52196 3072 52198
rect 3096 52196 3152 52198
rect 3176 52196 3232 52198
rect 3256 52196 3312 52198
rect 2356 51706 2412 51708
rect 2436 51706 2492 51708
rect 2516 51706 2572 51708
rect 2596 51706 2652 51708
rect 2356 51654 2402 51706
rect 2402 51654 2412 51706
rect 2436 51654 2466 51706
rect 2466 51654 2478 51706
rect 2478 51654 2492 51706
rect 2516 51654 2530 51706
rect 2530 51654 2542 51706
rect 2542 51654 2572 51706
rect 2596 51654 2606 51706
rect 2606 51654 2652 51706
rect 2356 51652 2412 51654
rect 2436 51652 2492 51654
rect 2516 51652 2572 51654
rect 2596 51652 2652 51654
rect 3016 51162 3072 51164
rect 3096 51162 3152 51164
rect 3176 51162 3232 51164
rect 3256 51162 3312 51164
rect 3016 51110 3062 51162
rect 3062 51110 3072 51162
rect 3096 51110 3126 51162
rect 3126 51110 3138 51162
rect 3138 51110 3152 51162
rect 3176 51110 3190 51162
rect 3190 51110 3202 51162
rect 3202 51110 3232 51162
rect 3256 51110 3266 51162
rect 3266 51110 3312 51162
rect 3016 51108 3072 51110
rect 3096 51108 3152 51110
rect 3176 51108 3232 51110
rect 3256 51108 3312 51110
rect 2356 50618 2412 50620
rect 2436 50618 2492 50620
rect 2516 50618 2572 50620
rect 2596 50618 2652 50620
rect 2356 50566 2402 50618
rect 2402 50566 2412 50618
rect 2436 50566 2466 50618
rect 2466 50566 2478 50618
rect 2478 50566 2492 50618
rect 2516 50566 2530 50618
rect 2530 50566 2542 50618
rect 2542 50566 2572 50618
rect 2596 50566 2606 50618
rect 2606 50566 2652 50618
rect 2356 50564 2412 50566
rect 2436 50564 2492 50566
rect 2516 50564 2572 50566
rect 2596 50564 2652 50566
rect 3016 50074 3072 50076
rect 3096 50074 3152 50076
rect 3176 50074 3232 50076
rect 3256 50074 3312 50076
rect 3016 50022 3062 50074
rect 3062 50022 3072 50074
rect 3096 50022 3126 50074
rect 3126 50022 3138 50074
rect 3138 50022 3152 50074
rect 3176 50022 3190 50074
rect 3190 50022 3202 50074
rect 3202 50022 3232 50074
rect 3256 50022 3266 50074
rect 3266 50022 3312 50074
rect 3016 50020 3072 50022
rect 3096 50020 3152 50022
rect 3176 50020 3232 50022
rect 3256 50020 3312 50022
rect 2356 49530 2412 49532
rect 2436 49530 2492 49532
rect 2516 49530 2572 49532
rect 2596 49530 2652 49532
rect 2356 49478 2402 49530
rect 2402 49478 2412 49530
rect 2436 49478 2466 49530
rect 2466 49478 2478 49530
rect 2478 49478 2492 49530
rect 2516 49478 2530 49530
rect 2530 49478 2542 49530
rect 2542 49478 2572 49530
rect 2596 49478 2606 49530
rect 2606 49478 2652 49530
rect 2356 49476 2412 49478
rect 2436 49476 2492 49478
rect 2516 49476 2572 49478
rect 2596 49476 2652 49478
rect 3016 48986 3072 48988
rect 3096 48986 3152 48988
rect 3176 48986 3232 48988
rect 3256 48986 3312 48988
rect 3016 48934 3062 48986
rect 3062 48934 3072 48986
rect 3096 48934 3126 48986
rect 3126 48934 3138 48986
rect 3138 48934 3152 48986
rect 3176 48934 3190 48986
rect 3190 48934 3202 48986
rect 3202 48934 3232 48986
rect 3256 48934 3266 48986
rect 3266 48934 3312 48986
rect 3016 48932 3072 48934
rect 3096 48932 3152 48934
rect 3176 48932 3232 48934
rect 3256 48932 3312 48934
rect 2356 48442 2412 48444
rect 2436 48442 2492 48444
rect 2516 48442 2572 48444
rect 2596 48442 2652 48444
rect 2356 48390 2402 48442
rect 2402 48390 2412 48442
rect 2436 48390 2466 48442
rect 2466 48390 2478 48442
rect 2478 48390 2492 48442
rect 2516 48390 2530 48442
rect 2530 48390 2542 48442
rect 2542 48390 2572 48442
rect 2596 48390 2606 48442
rect 2606 48390 2652 48442
rect 2356 48388 2412 48390
rect 2436 48388 2492 48390
rect 2516 48388 2572 48390
rect 2596 48388 2652 48390
rect 3016 47898 3072 47900
rect 3096 47898 3152 47900
rect 3176 47898 3232 47900
rect 3256 47898 3312 47900
rect 3016 47846 3062 47898
rect 3062 47846 3072 47898
rect 3096 47846 3126 47898
rect 3126 47846 3138 47898
rect 3138 47846 3152 47898
rect 3176 47846 3190 47898
rect 3190 47846 3202 47898
rect 3202 47846 3232 47898
rect 3256 47846 3266 47898
rect 3266 47846 3312 47898
rect 3016 47844 3072 47846
rect 3096 47844 3152 47846
rect 3176 47844 3232 47846
rect 3256 47844 3312 47846
rect 2356 47354 2412 47356
rect 2436 47354 2492 47356
rect 2516 47354 2572 47356
rect 2596 47354 2652 47356
rect 2356 47302 2402 47354
rect 2402 47302 2412 47354
rect 2436 47302 2466 47354
rect 2466 47302 2478 47354
rect 2478 47302 2492 47354
rect 2516 47302 2530 47354
rect 2530 47302 2542 47354
rect 2542 47302 2572 47354
rect 2596 47302 2606 47354
rect 2606 47302 2652 47354
rect 2356 47300 2412 47302
rect 2436 47300 2492 47302
rect 2516 47300 2572 47302
rect 2596 47300 2652 47302
rect 3016 46810 3072 46812
rect 3096 46810 3152 46812
rect 3176 46810 3232 46812
rect 3256 46810 3312 46812
rect 3016 46758 3062 46810
rect 3062 46758 3072 46810
rect 3096 46758 3126 46810
rect 3126 46758 3138 46810
rect 3138 46758 3152 46810
rect 3176 46758 3190 46810
rect 3190 46758 3202 46810
rect 3202 46758 3232 46810
rect 3256 46758 3266 46810
rect 3266 46758 3312 46810
rect 3016 46756 3072 46758
rect 3096 46756 3152 46758
rect 3176 46756 3232 46758
rect 3256 46756 3312 46758
rect 2356 46266 2412 46268
rect 2436 46266 2492 46268
rect 2516 46266 2572 46268
rect 2596 46266 2652 46268
rect 2356 46214 2402 46266
rect 2402 46214 2412 46266
rect 2436 46214 2466 46266
rect 2466 46214 2478 46266
rect 2478 46214 2492 46266
rect 2516 46214 2530 46266
rect 2530 46214 2542 46266
rect 2542 46214 2572 46266
rect 2596 46214 2606 46266
rect 2606 46214 2652 46266
rect 2356 46212 2412 46214
rect 2436 46212 2492 46214
rect 2516 46212 2572 46214
rect 2596 46212 2652 46214
rect 3016 45722 3072 45724
rect 3096 45722 3152 45724
rect 3176 45722 3232 45724
rect 3256 45722 3312 45724
rect 3016 45670 3062 45722
rect 3062 45670 3072 45722
rect 3096 45670 3126 45722
rect 3126 45670 3138 45722
rect 3138 45670 3152 45722
rect 3176 45670 3190 45722
rect 3190 45670 3202 45722
rect 3202 45670 3232 45722
rect 3256 45670 3266 45722
rect 3266 45670 3312 45722
rect 3016 45668 3072 45670
rect 3096 45668 3152 45670
rect 3176 45668 3232 45670
rect 3256 45668 3312 45670
rect 2356 45178 2412 45180
rect 2436 45178 2492 45180
rect 2516 45178 2572 45180
rect 2596 45178 2652 45180
rect 2356 45126 2402 45178
rect 2402 45126 2412 45178
rect 2436 45126 2466 45178
rect 2466 45126 2478 45178
rect 2478 45126 2492 45178
rect 2516 45126 2530 45178
rect 2530 45126 2542 45178
rect 2542 45126 2572 45178
rect 2596 45126 2606 45178
rect 2606 45126 2652 45178
rect 2356 45124 2412 45126
rect 2436 45124 2492 45126
rect 2516 45124 2572 45126
rect 2596 45124 2652 45126
rect 3016 44634 3072 44636
rect 3096 44634 3152 44636
rect 3176 44634 3232 44636
rect 3256 44634 3312 44636
rect 3016 44582 3062 44634
rect 3062 44582 3072 44634
rect 3096 44582 3126 44634
rect 3126 44582 3138 44634
rect 3138 44582 3152 44634
rect 3176 44582 3190 44634
rect 3190 44582 3202 44634
rect 3202 44582 3232 44634
rect 3256 44582 3266 44634
rect 3266 44582 3312 44634
rect 3016 44580 3072 44582
rect 3096 44580 3152 44582
rect 3176 44580 3232 44582
rect 3256 44580 3312 44582
rect 2356 44090 2412 44092
rect 2436 44090 2492 44092
rect 2516 44090 2572 44092
rect 2596 44090 2652 44092
rect 2356 44038 2402 44090
rect 2402 44038 2412 44090
rect 2436 44038 2466 44090
rect 2466 44038 2478 44090
rect 2478 44038 2492 44090
rect 2516 44038 2530 44090
rect 2530 44038 2542 44090
rect 2542 44038 2572 44090
rect 2596 44038 2606 44090
rect 2606 44038 2652 44090
rect 2356 44036 2412 44038
rect 2436 44036 2492 44038
rect 2516 44036 2572 44038
rect 2596 44036 2652 44038
rect 3016 43546 3072 43548
rect 3096 43546 3152 43548
rect 3176 43546 3232 43548
rect 3256 43546 3312 43548
rect 3016 43494 3062 43546
rect 3062 43494 3072 43546
rect 3096 43494 3126 43546
rect 3126 43494 3138 43546
rect 3138 43494 3152 43546
rect 3176 43494 3190 43546
rect 3190 43494 3202 43546
rect 3202 43494 3232 43546
rect 3256 43494 3266 43546
rect 3266 43494 3312 43546
rect 3016 43492 3072 43494
rect 3096 43492 3152 43494
rect 3176 43492 3232 43494
rect 3256 43492 3312 43494
rect 2356 43002 2412 43004
rect 2436 43002 2492 43004
rect 2516 43002 2572 43004
rect 2596 43002 2652 43004
rect 2356 42950 2402 43002
rect 2402 42950 2412 43002
rect 2436 42950 2466 43002
rect 2466 42950 2478 43002
rect 2478 42950 2492 43002
rect 2516 42950 2530 43002
rect 2530 42950 2542 43002
rect 2542 42950 2572 43002
rect 2596 42950 2606 43002
rect 2606 42950 2652 43002
rect 2356 42948 2412 42950
rect 2436 42948 2492 42950
rect 2516 42948 2572 42950
rect 2596 42948 2652 42950
rect 3016 42458 3072 42460
rect 3096 42458 3152 42460
rect 3176 42458 3232 42460
rect 3256 42458 3312 42460
rect 3016 42406 3062 42458
rect 3062 42406 3072 42458
rect 3096 42406 3126 42458
rect 3126 42406 3138 42458
rect 3138 42406 3152 42458
rect 3176 42406 3190 42458
rect 3190 42406 3202 42458
rect 3202 42406 3232 42458
rect 3256 42406 3266 42458
rect 3266 42406 3312 42458
rect 3016 42404 3072 42406
rect 3096 42404 3152 42406
rect 3176 42404 3232 42406
rect 3256 42404 3312 42406
rect 2356 41914 2412 41916
rect 2436 41914 2492 41916
rect 2516 41914 2572 41916
rect 2596 41914 2652 41916
rect 2356 41862 2402 41914
rect 2402 41862 2412 41914
rect 2436 41862 2466 41914
rect 2466 41862 2478 41914
rect 2478 41862 2492 41914
rect 2516 41862 2530 41914
rect 2530 41862 2542 41914
rect 2542 41862 2572 41914
rect 2596 41862 2606 41914
rect 2606 41862 2652 41914
rect 2356 41860 2412 41862
rect 2436 41860 2492 41862
rect 2516 41860 2572 41862
rect 2596 41860 2652 41862
rect 3016 41370 3072 41372
rect 3096 41370 3152 41372
rect 3176 41370 3232 41372
rect 3256 41370 3312 41372
rect 3016 41318 3062 41370
rect 3062 41318 3072 41370
rect 3096 41318 3126 41370
rect 3126 41318 3138 41370
rect 3138 41318 3152 41370
rect 3176 41318 3190 41370
rect 3190 41318 3202 41370
rect 3202 41318 3232 41370
rect 3256 41318 3266 41370
rect 3266 41318 3312 41370
rect 3016 41316 3072 41318
rect 3096 41316 3152 41318
rect 3176 41316 3232 41318
rect 3256 41316 3312 41318
rect 2356 40826 2412 40828
rect 2436 40826 2492 40828
rect 2516 40826 2572 40828
rect 2596 40826 2652 40828
rect 2356 40774 2402 40826
rect 2402 40774 2412 40826
rect 2436 40774 2466 40826
rect 2466 40774 2478 40826
rect 2478 40774 2492 40826
rect 2516 40774 2530 40826
rect 2530 40774 2542 40826
rect 2542 40774 2572 40826
rect 2596 40774 2606 40826
rect 2606 40774 2652 40826
rect 2356 40772 2412 40774
rect 2436 40772 2492 40774
rect 2516 40772 2572 40774
rect 2596 40772 2652 40774
rect 3016 40282 3072 40284
rect 3096 40282 3152 40284
rect 3176 40282 3232 40284
rect 3256 40282 3312 40284
rect 3016 40230 3062 40282
rect 3062 40230 3072 40282
rect 3096 40230 3126 40282
rect 3126 40230 3138 40282
rect 3138 40230 3152 40282
rect 3176 40230 3190 40282
rect 3190 40230 3202 40282
rect 3202 40230 3232 40282
rect 3256 40230 3266 40282
rect 3266 40230 3312 40282
rect 3016 40228 3072 40230
rect 3096 40228 3152 40230
rect 3176 40228 3232 40230
rect 3256 40228 3312 40230
rect 5630 40060 5632 40080
rect 5632 40060 5684 40080
rect 5684 40060 5686 40080
rect 5630 40024 5686 40060
rect 6182 41384 6238 41440
rect 6918 61240 6974 61296
rect 7356 77818 7412 77820
rect 7436 77818 7492 77820
rect 7516 77818 7572 77820
rect 7596 77818 7652 77820
rect 7356 77766 7402 77818
rect 7402 77766 7412 77818
rect 7436 77766 7466 77818
rect 7466 77766 7478 77818
rect 7478 77766 7492 77818
rect 7516 77766 7530 77818
rect 7530 77766 7542 77818
rect 7542 77766 7572 77818
rect 7596 77766 7606 77818
rect 7606 77766 7652 77818
rect 7356 77764 7412 77766
rect 7436 77764 7492 77766
rect 7516 77764 7572 77766
rect 7596 77764 7652 77766
rect 8016 77274 8072 77276
rect 8096 77274 8152 77276
rect 8176 77274 8232 77276
rect 8256 77274 8312 77276
rect 8016 77222 8062 77274
rect 8062 77222 8072 77274
rect 8096 77222 8126 77274
rect 8126 77222 8138 77274
rect 8138 77222 8152 77274
rect 8176 77222 8190 77274
rect 8190 77222 8202 77274
rect 8202 77222 8232 77274
rect 8256 77222 8266 77274
rect 8266 77222 8312 77274
rect 8016 77220 8072 77222
rect 8096 77220 8152 77222
rect 8176 77220 8232 77222
rect 8256 77220 8312 77222
rect 7356 76730 7412 76732
rect 7436 76730 7492 76732
rect 7516 76730 7572 76732
rect 7596 76730 7652 76732
rect 7356 76678 7402 76730
rect 7402 76678 7412 76730
rect 7436 76678 7466 76730
rect 7466 76678 7478 76730
rect 7478 76678 7492 76730
rect 7516 76678 7530 76730
rect 7530 76678 7542 76730
rect 7542 76678 7572 76730
rect 7596 76678 7606 76730
rect 7606 76678 7652 76730
rect 7356 76676 7412 76678
rect 7436 76676 7492 76678
rect 7516 76676 7572 76678
rect 7596 76676 7652 76678
rect 8016 76186 8072 76188
rect 8096 76186 8152 76188
rect 8176 76186 8232 76188
rect 8256 76186 8312 76188
rect 8016 76134 8062 76186
rect 8062 76134 8072 76186
rect 8096 76134 8126 76186
rect 8126 76134 8138 76186
rect 8138 76134 8152 76186
rect 8176 76134 8190 76186
rect 8190 76134 8202 76186
rect 8202 76134 8232 76186
rect 8256 76134 8266 76186
rect 8266 76134 8312 76186
rect 8016 76132 8072 76134
rect 8096 76132 8152 76134
rect 8176 76132 8232 76134
rect 8256 76132 8312 76134
rect 7356 75642 7412 75644
rect 7436 75642 7492 75644
rect 7516 75642 7572 75644
rect 7596 75642 7652 75644
rect 7356 75590 7402 75642
rect 7402 75590 7412 75642
rect 7436 75590 7466 75642
rect 7466 75590 7478 75642
rect 7478 75590 7492 75642
rect 7516 75590 7530 75642
rect 7530 75590 7542 75642
rect 7542 75590 7572 75642
rect 7596 75590 7606 75642
rect 7606 75590 7652 75642
rect 7356 75588 7412 75590
rect 7436 75588 7492 75590
rect 7516 75588 7572 75590
rect 7596 75588 7652 75590
rect 8016 75098 8072 75100
rect 8096 75098 8152 75100
rect 8176 75098 8232 75100
rect 8256 75098 8312 75100
rect 8016 75046 8062 75098
rect 8062 75046 8072 75098
rect 8096 75046 8126 75098
rect 8126 75046 8138 75098
rect 8138 75046 8152 75098
rect 8176 75046 8190 75098
rect 8190 75046 8202 75098
rect 8202 75046 8232 75098
rect 8256 75046 8266 75098
rect 8266 75046 8312 75098
rect 8016 75044 8072 75046
rect 8096 75044 8152 75046
rect 8176 75044 8232 75046
rect 8256 75044 8312 75046
rect 7356 74554 7412 74556
rect 7436 74554 7492 74556
rect 7516 74554 7572 74556
rect 7596 74554 7652 74556
rect 7356 74502 7402 74554
rect 7402 74502 7412 74554
rect 7436 74502 7466 74554
rect 7466 74502 7478 74554
rect 7478 74502 7492 74554
rect 7516 74502 7530 74554
rect 7530 74502 7542 74554
rect 7542 74502 7572 74554
rect 7596 74502 7606 74554
rect 7606 74502 7652 74554
rect 7356 74500 7412 74502
rect 7436 74500 7492 74502
rect 7516 74500 7572 74502
rect 7596 74500 7652 74502
rect 8016 74010 8072 74012
rect 8096 74010 8152 74012
rect 8176 74010 8232 74012
rect 8256 74010 8312 74012
rect 8016 73958 8062 74010
rect 8062 73958 8072 74010
rect 8096 73958 8126 74010
rect 8126 73958 8138 74010
rect 8138 73958 8152 74010
rect 8176 73958 8190 74010
rect 8190 73958 8202 74010
rect 8202 73958 8232 74010
rect 8256 73958 8266 74010
rect 8266 73958 8312 74010
rect 8016 73956 8072 73958
rect 8096 73956 8152 73958
rect 8176 73956 8232 73958
rect 8256 73956 8312 73958
rect 7356 73466 7412 73468
rect 7436 73466 7492 73468
rect 7516 73466 7572 73468
rect 7596 73466 7652 73468
rect 7356 73414 7402 73466
rect 7402 73414 7412 73466
rect 7436 73414 7466 73466
rect 7466 73414 7478 73466
rect 7478 73414 7492 73466
rect 7516 73414 7530 73466
rect 7530 73414 7542 73466
rect 7542 73414 7572 73466
rect 7596 73414 7606 73466
rect 7606 73414 7652 73466
rect 7356 73412 7412 73414
rect 7436 73412 7492 73414
rect 7516 73412 7572 73414
rect 7596 73412 7652 73414
rect 7356 72378 7412 72380
rect 7436 72378 7492 72380
rect 7516 72378 7572 72380
rect 7596 72378 7652 72380
rect 7356 72326 7402 72378
rect 7402 72326 7412 72378
rect 7436 72326 7466 72378
rect 7466 72326 7478 72378
rect 7478 72326 7492 72378
rect 7516 72326 7530 72378
rect 7530 72326 7542 72378
rect 7542 72326 7572 72378
rect 7596 72326 7606 72378
rect 7606 72326 7652 72378
rect 7356 72324 7412 72326
rect 7436 72324 7492 72326
rect 7516 72324 7572 72326
rect 7596 72324 7652 72326
rect 8390 73208 8446 73264
rect 8016 72922 8072 72924
rect 8096 72922 8152 72924
rect 8176 72922 8232 72924
rect 8256 72922 8312 72924
rect 8016 72870 8062 72922
rect 8062 72870 8072 72922
rect 8096 72870 8126 72922
rect 8126 72870 8138 72922
rect 8138 72870 8152 72922
rect 8176 72870 8190 72922
rect 8190 72870 8202 72922
rect 8202 72870 8232 72922
rect 8256 72870 8266 72922
rect 8266 72870 8312 72922
rect 8016 72868 8072 72870
rect 8096 72868 8152 72870
rect 8176 72868 8232 72870
rect 8256 72868 8312 72870
rect 8482 71848 8538 71904
rect 8016 71834 8072 71836
rect 8096 71834 8152 71836
rect 8176 71834 8232 71836
rect 8256 71834 8312 71836
rect 8016 71782 8062 71834
rect 8062 71782 8072 71834
rect 8096 71782 8126 71834
rect 8126 71782 8138 71834
rect 8138 71782 8152 71834
rect 8176 71782 8190 71834
rect 8190 71782 8202 71834
rect 8202 71782 8232 71834
rect 8256 71782 8266 71834
rect 8266 71782 8312 71834
rect 8016 71780 8072 71782
rect 8096 71780 8152 71782
rect 8176 71780 8232 71782
rect 8256 71780 8312 71782
rect 7356 71290 7412 71292
rect 7436 71290 7492 71292
rect 7516 71290 7572 71292
rect 7596 71290 7652 71292
rect 7356 71238 7402 71290
rect 7402 71238 7412 71290
rect 7436 71238 7466 71290
rect 7466 71238 7478 71290
rect 7478 71238 7492 71290
rect 7516 71238 7530 71290
rect 7530 71238 7542 71290
rect 7542 71238 7572 71290
rect 7596 71238 7606 71290
rect 7606 71238 7652 71290
rect 7356 71236 7412 71238
rect 7436 71236 7492 71238
rect 7516 71236 7572 71238
rect 7596 71236 7652 71238
rect 7356 70202 7412 70204
rect 7436 70202 7492 70204
rect 7516 70202 7572 70204
rect 7596 70202 7652 70204
rect 7356 70150 7402 70202
rect 7402 70150 7412 70202
rect 7436 70150 7466 70202
rect 7466 70150 7478 70202
rect 7478 70150 7492 70202
rect 7516 70150 7530 70202
rect 7530 70150 7542 70202
rect 7542 70150 7572 70202
rect 7596 70150 7606 70202
rect 7606 70150 7652 70202
rect 7356 70148 7412 70150
rect 7436 70148 7492 70150
rect 7516 70148 7572 70150
rect 7596 70148 7652 70150
rect 8016 70746 8072 70748
rect 8096 70746 8152 70748
rect 8176 70746 8232 70748
rect 8256 70746 8312 70748
rect 8016 70694 8062 70746
rect 8062 70694 8072 70746
rect 8096 70694 8126 70746
rect 8126 70694 8138 70746
rect 8138 70694 8152 70746
rect 8176 70694 8190 70746
rect 8190 70694 8202 70746
rect 8202 70694 8232 70746
rect 8256 70694 8266 70746
rect 8266 70694 8312 70746
rect 8016 70692 8072 70694
rect 8096 70692 8152 70694
rect 8176 70692 8232 70694
rect 8256 70692 8312 70694
rect 8390 70488 8446 70544
rect 8016 69658 8072 69660
rect 8096 69658 8152 69660
rect 8176 69658 8232 69660
rect 8256 69658 8312 69660
rect 8016 69606 8062 69658
rect 8062 69606 8072 69658
rect 8096 69606 8126 69658
rect 8126 69606 8138 69658
rect 8138 69606 8152 69658
rect 8176 69606 8190 69658
rect 8190 69606 8202 69658
rect 8202 69606 8232 69658
rect 8256 69606 8266 69658
rect 8266 69606 8312 69658
rect 8016 69604 8072 69606
rect 8096 69604 8152 69606
rect 8176 69604 8232 69606
rect 8256 69604 8312 69606
rect 7356 69114 7412 69116
rect 7436 69114 7492 69116
rect 7516 69114 7572 69116
rect 7596 69114 7652 69116
rect 7356 69062 7402 69114
rect 7402 69062 7412 69114
rect 7436 69062 7466 69114
rect 7466 69062 7478 69114
rect 7478 69062 7492 69114
rect 7516 69062 7530 69114
rect 7530 69062 7542 69114
rect 7542 69062 7572 69114
rect 7596 69062 7606 69114
rect 7606 69062 7652 69114
rect 7356 69060 7412 69062
rect 7436 69060 7492 69062
rect 7516 69060 7572 69062
rect 7596 69060 7652 69062
rect 8390 69164 8392 69184
rect 8392 69164 8444 69184
rect 8444 69164 8446 69184
rect 8390 69128 8446 69164
rect 8016 68570 8072 68572
rect 8096 68570 8152 68572
rect 8176 68570 8232 68572
rect 8256 68570 8312 68572
rect 8016 68518 8062 68570
rect 8062 68518 8072 68570
rect 8096 68518 8126 68570
rect 8126 68518 8138 68570
rect 8138 68518 8152 68570
rect 8176 68518 8190 68570
rect 8190 68518 8202 68570
rect 8202 68518 8232 68570
rect 8256 68518 8266 68570
rect 8266 68518 8312 68570
rect 8016 68516 8072 68518
rect 8096 68516 8152 68518
rect 8176 68516 8232 68518
rect 8256 68516 8312 68518
rect 7356 68026 7412 68028
rect 7436 68026 7492 68028
rect 7516 68026 7572 68028
rect 7596 68026 7652 68028
rect 7356 67974 7402 68026
rect 7402 67974 7412 68026
rect 7436 67974 7466 68026
rect 7466 67974 7478 68026
rect 7478 67974 7492 68026
rect 7516 67974 7530 68026
rect 7530 67974 7542 68026
rect 7542 67974 7572 68026
rect 7596 67974 7606 68026
rect 7606 67974 7652 68026
rect 7356 67972 7412 67974
rect 7436 67972 7492 67974
rect 7516 67972 7572 67974
rect 7596 67972 7652 67974
rect 7356 66938 7412 66940
rect 7436 66938 7492 66940
rect 7516 66938 7572 66940
rect 7596 66938 7652 66940
rect 7356 66886 7402 66938
rect 7402 66886 7412 66938
rect 7436 66886 7466 66938
rect 7466 66886 7478 66938
rect 7478 66886 7492 66938
rect 7516 66886 7530 66938
rect 7530 66886 7542 66938
rect 7542 66886 7572 66938
rect 7596 66886 7606 66938
rect 7606 66886 7652 66938
rect 7356 66884 7412 66886
rect 7436 66884 7492 66886
rect 7516 66884 7572 66886
rect 7596 66884 7652 66886
rect 7356 65850 7412 65852
rect 7436 65850 7492 65852
rect 7516 65850 7572 65852
rect 7596 65850 7652 65852
rect 7356 65798 7402 65850
rect 7402 65798 7412 65850
rect 7436 65798 7466 65850
rect 7466 65798 7478 65850
rect 7478 65798 7492 65850
rect 7516 65798 7530 65850
rect 7530 65798 7542 65850
rect 7542 65798 7572 65850
rect 7596 65798 7606 65850
rect 7606 65798 7652 65850
rect 7356 65796 7412 65798
rect 7436 65796 7492 65798
rect 7516 65796 7572 65798
rect 7596 65796 7652 65798
rect 8390 67768 8446 67824
rect 8016 67482 8072 67484
rect 8096 67482 8152 67484
rect 8176 67482 8232 67484
rect 8256 67482 8312 67484
rect 8016 67430 8062 67482
rect 8062 67430 8072 67482
rect 8096 67430 8126 67482
rect 8126 67430 8138 67482
rect 8138 67430 8152 67482
rect 8176 67430 8190 67482
rect 8190 67430 8202 67482
rect 8202 67430 8232 67482
rect 8256 67430 8266 67482
rect 8266 67430 8312 67482
rect 8016 67428 8072 67430
rect 8096 67428 8152 67430
rect 8176 67428 8232 67430
rect 8256 67428 8312 67430
rect 8390 66408 8446 66464
rect 8016 66394 8072 66396
rect 8096 66394 8152 66396
rect 8176 66394 8232 66396
rect 8256 66394 8312 66396
rect 8016 66342 8062 66394
rect 8062 66342 8072 66394
rect 8096 66342 8126 66394
rect 8126 66342 8138 66394
rect 8138 66342 8152 66394
rect 8176 66342 8190 66394
rect 8190 66342 8202 66394
rect 8202 66342 8232 66394
rect 8256 66342 8266 66394
rect 8266 66342 8312 66394
rect 8016 66340 8072 66342
rect 8096 66340 8152 66342
rect 8176 66340 8232 66342
rect 8256 66340 8312 66342
rect 7356 64762 7412 64764
rect 7436 64762 7492 64764
rect 7516 64762 7572 64764
rect 7596 64762 7652 64764
rect 7356 64710 7402 64762
rect 7402 64710 7412 64762
rect 7436 64710 7466 64762
rect 7466 64710 7478 64762
rect 7478 64710 7492 64762
rect 7516 64710 7530 64762
rect 7530 64710 7542 64762
rect 7542 64710 7572 64762
rect 7596 64710 7606 64762
rect 7606 64710 7652 64762
rect 7356 64708 7412 64710
rect 7436 64708 7492 64710
rect 7516 64708 7572 64710
rect 7596 64708 7652 64710
rect 7356 63674 7412 63676
rect 7436 63674 7492 63676
rect 7516 63674 7572 63676
rect 7596 63674 7652 63676
rect 7356 63622 7402 63674
rect 7402 63622 7412 63674
rect 7436 63622 7466 63674
rect 7466 63622 7478 63674
rect 7478 63622 7492 63674
rect 7516 63622 7530 63674
rect 7530 63622 7542 63674
rect 7542 63622 7572 63674
rect 7596 63622 7606 63674
rect 7606 63622 7652 63674
rect 7356 63620 7412 63622
rect 7436 63620 7492 63622
rect 7516 63620 7572 63622
rect 7596 63620 7652 63622
rect 7356 62586 7412 62588
rect 7436 62586 7492 62588
rect 7516 62586 7572 62588
rect 7596 62586 7652 62588
rect 7356 62534 7402 62586
rect 7402 62534 7412 62586
rect 7436 62534 7466 62586
rect 7466 62534 7478 62586
rect 7478 62534 7492 62586
rect 7516 62534 7530 62586
rect 7530 62534 7542 62586
rect 7542 62534 7572 62586
rect 7596 62534 7606 62586
rect 7606 62534 7652 62586
rect 7356 62532 7412 62534
rect 7436 62532 7492 62534
rect 7516 62532 7572 62534
rect 7596 62532 7652 62534
rect 7356 61498 7412 61500
rect 7436 61498 7492 61500
rect 7516 61498 7572 61500
rect 7596 61498 7652 61500
rect 7356 61446 7402 61498
rect 7402 61446 7412 61498
rect 7436 61446 7466 61498
rect 7466 61446 7478 61498
rect 7478 61446 7492 61498
rect 7516 61446 7530 61498
rect 7530 61446 7542 61498
rect 7542 61446 7572 61498
rect 7596 61446 7606 61498
rect 7606 61446 7652 61498
rect 7356 61444 7412 61446
rect 7436 61444 7492 61446
rect 7516 61444 7572 61446
rect 7596 61444 7652 61446
rect 8016 65306 8072 65308
rect 8096 65306 8152 65308
rect 8176 65306 8232 65308
rect 8256 65306 8312 65308
rect 8016 65254 8062 65306
rect 8062 65254 8072 65306
rect 8096 65254 8126 65306
rect 8126 65254 8138 65306
rect 8138 65254 8152 65306
rect 8176 65254 8190 65306
rect 8190 65254 8202 65306
rect 8202 65254 8232 65306
rect 8256 65254 8266 65306
rect 8266 65254 8312 65306
rect 8016 65252 8072 65254
rect 8096 65252 8152 65254
rect 8176 65252 8232 65254
rect 8256 65252 8312 65254
rect 8390 65048 8446 65104
rect 8016 64218 8072 64220
rect 8096 64218 8152 64220
rect 8176 64218 8232 64220
rect 8256 64218 8312 64220
rect 8016 64166 8062 64218
rect 8062 64166 8072 64218
rect 8096 64166 8126 64218
rect 8126 64166 8138 64218
rect 8138 64166 8152 64218
rect 8176 64166 8190 64218
rect 8190 64166 8202 64218
rect 8202 64166 8232 64218
rect 8256 64166 8266 64218
rect 8266 64166 8312 64218
rect 8016 64164 8072 64166
rect 8096 64164 8152 64166
rect 8176 64164 8232 64166
rect 8256 64164 8312 64166
rect 8482 63688 8538 63744
rect 8016 63130 8072 63132
rect 8096 63130 8152 63132
rect 8176 63130 8232 63132
rect 8256 63130 8312 63132
rect 8016 63078 8062 63130
rect 8062 63078 8072 63130
rect 8096 63078 8126 63130
rect 8126 63078 8138 63130
rect 8138 63078 8152 63130
rect 8176 63078 8190 63130
rect 8190 63078 8202 63130
rect 8202 63078 8232 63130
rect 8256 63078 8266 63130
rect 8266 63078 8312 63130
rect 8016 63076 8072 63078
rect 8096 63076 8152 63078
rect 8176 63076 8232 63078
rect 8256 63076 8312 63078
rect 8390 62328 8446 62384
rect 8016 62042 8072 62044
rect 8096 62042 8152 62044
rect 8176 62042 8232 62044
rect 8256 62042 8312 62044
rect 8016 61990 8062 62042
rect 8062 61990 8072 62042
rect 8096 61990 8126 62042
rect 8126 61990 8138 62042
rect 8138 61990 8152 62042
rect 8176 61990 8190 62042
rect 8190 61990 8202 62042
rect 8202 61990 8232 62042
rect 8256 61990 8266 62042
rect 8266 61990 8312 62042
rect 8016 61988 8072 61990
rect 8096 61988 8152 61990
rect 8176 61988 8232 61990
rect 8256 61988 8312 61990
rect 7838 60560 7894 60616
rect 7356 60410 7412 60412
rect 7436 60410 7492 60412
rect 7516 60410 7572 60412
rect 7596 60410 7652 60412
rect 7356 60358 7402 60410
rect 7402 60358 7412 60410
rect 7436 60358 7466 60410
rect 7466 60358 7478 60410
rect 7478 60358 7492 60410
rect 7516 60358 7530 60410
rect 7530 60358 7542 60410
rect 7542 60358 7572 60410
rect 7596 60358 7606 60410
rect 7606 60358 7652 60410
rect 7356 60356 7412 60358
rect 7436 60356 7492 60358
rect 7516 60356 7572 60358
rect 7596 60356 7652 60358
rect 7356 59322 7412 59324
rect 7436 59322 7492 59324
rect 7516 59322 7572 59324
rect 7596 59322 7652 59324
rect 7356 59270 7402 59322
rect 7402 59270 7412 59322
rect 7436 59270 7466 59322
rect 7466 59270 7478 59322
rect 7478 59270 7492 59322
rect 7516 59270 7530 59322
rect 7530 59270 7542 59322
rect 7542 59270 7572 59322
rect 7596 59270 7606 59322
rect 7606 59270 7652 59322
rect 7356 59268 7412 59270
rect 7436 59268 7492 59270
rect 7516 59268 7572 59270
rect 7596 59268 7652 59270
rect 7356 58234 7412 58236
rect 7436 58234 7492 58236
rect 7516 58234 7572 58236
rect 7596 58234 7652 58236
rect 7356 58182 7402 58234
rect 7402 58182 7412 58234
rect 7436 58182 7466 58234
rect 7466 58182 7478 58234
rect 7478 58182 7492 58234
rect 7516 58182 7530 58234
rect 7530 58182 7542 58234
rect 7542 58182 7572 58234
rect 7596 58182 7606 58234
rect 7606 58182 7652 58234
rect 7356 58180 7412 58182
rect 7436 58180 7492 58182
rect 7516 58180 7572 58182
rect 7596 58180 7652 58182
rect 7356 57146 7412 57148
rect 7436 57146 7492 57148
rect 7516 57146 7572 57148
rect 7596 57146 7652 57148
rect 7356 57094 7402 57146
rect 7402 57094 7412 57146
rect 7436 57094 7466 57146
rect 7466 57094 7478 57146
rect 7478 57094 7492 57146
rect 7516 57094 7530 57146
rect 7530 57094 7542 57146
rect 7542 57094 7572 57146
rect 7596 57094 7606 57146
rect 7606 57094 7652 57146
rect 7356 57092 7412 57094
rect 7436 57092 7492 57094
rect 7516 57092 7572 57094
rect 7596 57092 7652 57094
rect 7356 56058 7412 56060
rect 7436 56058 7492 56060
rect 7516 56058 7572 56060
rect 7596 56058 7652 56060
rect 7356 56006 7402 56058
rect 7402 56006 7412 56058
rect 7436 56006 7466 56058
rect 7466 56006 7478 56058
rect 7478 56006 7492 56058
rect 7516 56006 7530 56058
rect 7530 56006 7542 56058
rect 7542 56006 7572 56058
rect 7596 56006 7606 56058
rect 7606 56006 7652 56058
rect 7356 56004 7412 56006
rect 7436 56004 7492 56006
rect 7516 56004 7572 56006
rect 7596 56004 7652 56006
rect 7356 54970 7412 54972
rect 7436 54970 7492 54972
rect 7516 54970 7572 54972
rect 7596 54970 7652 54972
rect 7356 54918 7402 54970
rect 7402 54918 7412 54970
rect 7436 54918 7466 54970
rect 7466 54918 7478 54970
rect 7478 54918 7492 54970
rect 7516 54918 7530 54970
rect 7530 54918 7542 54970
rect 7542 54918 7572 54970
rect 7596 54918 7606 54970
rect 7606 54918 7652 54970
rect 7356 54916 7412 54918
rect 7436 54916 7492 54918
rect 7516 54916 7572 54918
rect 7596 54916 7652 54918
rect 7356 53882 7412 53884
rect 7436 53882 7492 53884
rect 7516 53882 7572 53884
rect 7596 53882 7652 53884
rect 7356 53830 7402 53882
rect 7402 53830 7412 53882
rect 7436 53830 7466 53882
rect 7466 53830 7478 53882
rect 7478 53830 7492 53882
rect 7516 53830 7530 53882
rect 7530 53830 7542 53882
rect 7542 53830 7572 53882
rect 7596 53830 7606 53882
rect 7606 53830 7652 53882
rect 7356 53828 7412 53830
rect 7436 53828 7492 53830
rect 7516 53828 7572 53830
rect 7596 53828 7652 53830
rect 7356 52794 7412 52796
rect 7436 52794 7492 52796
rect 7516 52794 7572 52796
rect 7596 52794 7652 52796
rect 7356 52742 7402 52794
rect 7402 52742 7412 52794
rect 7436 52742 7466 52794
rect 7466 52742 7478 52794
rect 7478 52742 7492 52794
rect 7516 52742 7530 52794
rect 7530 52742 7542 52794
rect 7542 52742 7572 52794
rect 7596 52742 7606 52794
rect 7606 52742 7652 52794
rect 7356 52740 7412 52742
rect 7436 52740 7492 52742
rect 7516 52740 7572 52742
rect 7596 52740 7652 52742
rect 7356 51706 7412 51708
rect 7436 51706 7492 51708
rect 7516 51706 7572 51708
rect 7596 51706 7652 51708
rect 7356 51654 7402 51706
rect 7402 51654 7412 51706
rect 7436 51654 7466 51706
rect 7466 51654 7478 51706
rect 7478 51654 7492 51706
rect 7516 51654 7530 51706
rect 7530 51654 7542 51706
rect 7542 51654 7572 51706
rect 7596 51654 7606 51706
rect 7606 51654 7652 51706
rect 7356 51652 7412 51654
rect 7436 51652 7492 51654
rect 7516 51652 7572 51654
rect 7596 51652 7652 51654
rect 8390 61004 8392 61024
rect 8392 61004 8444 61024
rect 8444 61004 8446 61024
rect 8390 60968 8446 61004
rect 8016 60954 8072 60956
rect 8096 60954 8152 60956
rect 8176 60954 8232 60956
rect 8256 60954 8312 60956
rect 8016 60902 8062 60954
rect 8062 60902 8072 60954
rect 8096 60902 8126 60954
rect 8126 60902 8138 60954
rect 8138 60902 8152 60954
rect 8176 60902 8190 60954
rect 8190 60902 8202 60954
rect 8202 60902 8232 60954
rect 8256 60902 8266 60954
rect 8266 60902 8312 60954
rect 8016 60900 8072 60902
rect 8096 60900 8152 60902
rect 8176 60900 8232 60902
rect 8256 60900 8312 60902
rect 8016 59866 8072 59868
rect 8096 59866 8152 59868
rect 8176 59866 8232 59868
rect 8256 59866 8312 59868
rect 8016 59814 8062 59866
rect 8062 59814 8072 59866
rect 8096 59814 8126 59866
rect 8126 59814 8138 59866
rect 8138 59814 8152 59866
rect 8176 59814 8190 59866
rect 8190 59814 8202 59866
rect 8202 59814 8232 59866
rect 8256 59814 8266 59866
rect 8266 59814 8312 59866
rect 8016 59812 8072 59814
rect 8096 59812 8152 59814
rect 8176 59812 8232 59814
rect 8256 59812 8312 59814
rect 8390 59608 8446 59664
rect 8016 58778 8072 58780
rect 8096 58778 8152 58780
rect 8176 58778 8232 58780
rect 8256 58778 8312 58780
rect 8016 58726 8062 58778
rect 8062 58726 8072 58778
rect 8096 58726 8126 58778
rect 8126 58726 8138 58778
rect 8138 58726 8152 58778
rect 8176 58726 8190 58778
rect 8190 58726 8202 58778
rect 8202 58726 8232 58778
rect 8256 58726 8266 58778
rect 8266 58726 8312 58778
rect 8016 58724 8072 58726
rect 8096 58724 8152 58726
rect 8176 58724 8232 58726
rect 8256 58724 8312 58726
rect 8482 58248 8538 58304
rect 8016 57690 8072 57692
rect 8096 57690 8152 57692
rect 8176 57690 8232 57692
rect 8256 57690 8312 57692
rect 8016 57638 8062 57690
rect 8062 57638 8072 57690
rect 8096 57638 8126 57690
rect 8126 57638 8138 57690
rect 8138 57638 8152 57690
rect 8176 57638 8190 57690
rect 8190 57638 8202 57690
rect 8202 57638 8232 57690
rect 8256 57638 8266 57690
rect 8266 57638 8312 57690
rect 8016 57636 8072 57638
rect 8096 57636 8152 57638
rect 8176 57636 8232 57638
rect 8256 57636 8312 57638
rect 8574 56888 8630 56944
rect 8016 56602 8072 56604
rect 8096 56602 8152 56604
rect 8176 56602 8232 56604
rect 8256 56602 8312 56604
rect 8016 56550 8062 56602
rect 8062 56550 8072 56602
rect 8096 56550 8126 56602
rect 8126 56550 8138 56602
rect 8138 56550 8152 56602
rect 8176 56550 8190 56602
rect 8190 56550 8202 56602
rect 8202 56550 8232 56602
rect 8256 56550 8266 56602
rect 8266 56550 8312 56602
rect 8016 56548 8072 56550
rect 8096 56548 8152 56550
rect 8176 56548 8232 56550
rect 8256 56548 8312 56550
rect 8016 55514 8072 55516
rect 8096 55514 8152 55516
rect 8176 55514 8232 55516
rect 8256 55514 8312 55516
rect 8016 55462 8062 55514
rect 8062 55462 8072 55514
rect 8096 55462 8126 55514
rect 8126 55462 8138 55514
rect 8138 55462 8152 55514
rect 8176 55462 8190 55514
rect 8190 55462 8202 55514
rect 8202 55462 8232 55514
rect 8256 55462 8266 55514
rect 8266 55462 8312 55514
rect 8016 55460 8072 55462
rect 8096 55460 8152 55462
rect 8176 55460 8232 55462
rect 8256 55460 8312 55462
rect 8206 55256 8262 55312
rect 8016 54426 8072 54428
rect 8096 54426 8152 54428
rect 8176 54426 8232 54428
rect 8256 54426 8312 54428
rect 8016 54374 8062 54426
rect 8062 54374 8072 54426
rect 8096 54374 8126 54426
rect 8126 54374 8138 54426
rect 8138 54374 8152 54426
rect 8176 54374 8190 54426
rect 8190 54374 8202 54426
rect 8202 54374 8232 54426
rect 8256 54374 8266 54426
rect 8266 54374 8312 54426
rect 8016 54372 8072 54374
rect 8096 54372 8152 54374
rect 8176 54372 8232 54374
rect 8256 54372 8312 54374
rect 8390 54168 8446 54224
rect 8016 53338 8072 53340
rect 8096 53338 8152 53340
rect 8176 53338 8232 53340
rect 8256 53338 8312 53340
rect 8016 53286 8062 53338
rect 8062 53286 8072 53338
rect 8096 53286 8126 53338
rect 8126 53286 8138 53338
rect 8138 53286 8152 53338
rect 8176 53286 8190 53338
rect 8190 53286 8202 53338
rect 8202 53286 8232 53338
rect 8256 53286 8266 53338
rect 8266 53286 8312 53338
rect 8016 53284 8072 53286
rect 8096 53284 8152 53286
rect 8176 53284 8232 53286
rect 8256 53284 8312 53286
rect 8390 52808 8446 52864
rect 8016 52250 8072 52252
rect 8096 52250 8152 52252
rect 8176 52250 8232 52252
rect 8256 52250 8312 52252
rect 8016 52198 8062 52250
rect 8062 52198 8072 52250
rect 8096 52198 8126 52250
rect 8126 52198 8138 52250
rect 8138 52198 8152 52250
rect 8176 52198 8190 52250
rect 8190 52198 8202 52250
rect 8202 52198 8232 52250
rect 8256 52198 8266 52250
rect 8266 52198 8312 52250
rect 8016 52196 8072 52198
rect 8096 52196 8152 52198
rect 8176 52196 8232 52198
rect 8256 52196 8312 52198
rect 8390 51448 8446 51504
rect 8016 51162 8072 51164
rect 8096 51162 8152 51164
rect 8176 51162 8232 51164
rect 8256 51162 8312 51164
rect 8016 51110 8062 51162
rect 8062 51110 8072 51162
rect 8096 51110 8126 51162
rect 8126 51110 8138 51162
rect 8138 51110 8152 51162
rect 8176 51110 8190 51162
rect 8190 51110 8202 51162
rect 8202 51110 8232 51162
rect 8256 51110 8266 51162
rect 8266 51110 8312 51162
rect 8016 51108 8072 51110
rect 8096 51108 8152 51110
rect 8176 51108 8232 51110
rect 8256 51108 8312 51110
rect 7356 50618 7412 50620
rect 7436 50618 7492 50620
rect 7516 50618 7572 50620
rect 7596 50618 7652 50620
rect 7356 50566 7402 50618
rect 7402 50566 7412 50618
rect 7436 50566 7466 50618
rect 7466 50566 7478 50618
rect 7478 50566 7492 50618
rect 7516 50566 7530 50618
rect 7530 50566 7542 50618
rect 7542 50566 7572 50618
rect 7596 50566 7606 50618
rect 7606 50566 7652 50618
rect 7356 50564 7412 50566
rect 7436 50564 7492 50566
rect 7516 50564 7572 50566
rect 7596 50564 7652 50566
rect 7356 49530 7412 49532
rect 7436 49530 7492 49532
rect 7516 49530 7572 49532
rect 7596 49530 7652 49532
rect 7356 49478 7402 49530
rect 7402 49478 7412 49530
rect 7436 49478 7466 49530
rect 7466 49478 7478 49530
rect 7478 49478 7492 49530
rect 7516 49478 7530 49530
rect 7530 49478 7542 49530
rect 7542 49478 7572 49530
rect 7596 49478 7606 49530
rect 7606 49478 7652 49530
rect 7356 49476 7412 49478
rect 7436 49476 7492 49478
rect 7516 49476 7572 49478
rect 7596 49476 7652 49478
rect 7356 48442 7412 48444
rect 7436 48442 7492 48444
rect 7516 48442 7572 48444
rect 7596 48442 7652 48444
rect 7356 48390 7402 48442
rect 7402 48390 7412 48442
rect 7436 48390 7466 48442
rect 7466 48390 7478 48442
rect 7478 48390 7492 48442
rect 7516 48390 7530 48442
rect 7530 48390 7542 48442
rect 7542 48390 7572 48442
rect 7596 48390 7606 48442
rect 7606 48390 7652 48442
rect 7356 48388 7412 48390
rect 7436 48388 7492 48390
rect 7516 48388 7572 48390
rect 7596 48388 7652 48390
rect 8390 50088 8446 50144
rect 8016 50074 8072 50076
rect 8096 50074 8152 50076
rect 8176 50074 8232 50076
rect 8256 50074 8312 50076
rect 8016 50022 8062 50074
rect 8062 50022 8072 50074
rect 8096 50022 8126 50074
rect 8126 50022 8138 50074
rect 8138 50022 8152 50074
rect 8176 50022 8190 50074
rect 8190 50022 8202 50074
rect 8202 50022 8232 50074
rect 8256 50022 8266 50074
rect 8266 50022 8312 50074
rect 8016 50020 8072 50022
rect 8096 50020 8152 50022
rect 8176 50020 8232 50022
rect 8256 50020 8312 50022
rect 8016 48986 8072 48988
rect 8096 48986 8152 48988
rect 8176 48986 8232 48988
rect 8256 48986 8312 48988
rect 8016 48934 8062 48986
rect 8062 48934 8072 48986
rect 8096 48934 8126 48986
rect 8126 48934 8138 48986
rect 8138 48934 8152 48986
rect 8176 48934 8190 48986
rect 8190 48934 8202 48986
rect 8202 48934 8232 48986
rect 8256 48934 8266 48986
rect 8266 48934 8312 48986
rect 8016 48932 8072 48934
rect 8096 48932 8152 48934
rect 8176 48932 8232 48934
rect 8256 48932 8312 48934
rect 8390 48728 8446 48784
rect 7356 47354 7412 47356
rect 7436 47354 7492 47356
rect 7516 47354 7572 47356
rect 7596 47354 7652 47356
rect 7356 47302 7402 47354
rect 7402 47302 7412 47354
rect 7436 47302 7466 47354
rect 7466 47302 7478 47354
rect 7478 47302 7492 47354
rect 7516 47302 7530 47354
rect 7530 47302 7542 47354
rect 7542 47302 7572 47354
rect 7596 47302 7606 47354
rect 7606 47302 7652 47354
rect 7356 47300 7412 47302
rect 7436 47300 7492 47302
rect 7516 47300 7572 47302
rect 7596 47300 7652 47302
rect 7356 46266 7412 46268
rect 7436 46266 7492 46268
rect 7516 46266 7572 46268
rect 7596 46266 7652 46268
rect 7356 46214 7402 46266
rect 7402 46214 7412 46266
rect 7436 46214 7466 46266
rect 7466 46214 7478 46266
rect 7478 46214 7492 46266
rect 7516 46214 7530 46266
rect 7530 46214 7542 46266
rect 7542 46214 7572 46266
rect 7596 46214 7606 46266
rect 7606 46214 7652 46266
rect 7356 46212 7412 46214
rect 7436 46212 7492 46214
rect 7516 46212 7572 46214
rect 7596 46212 7652 46214
rect 2356 39738 2412 39740
rect 2436 39738 2492 39740
rect 2516 39738 2572 39740
rect 2596 39738 2652 39740
rect 2356 39686 2402 39738
rect 2402 39686 2412 39738
rect 2436 39686 2466 39738
rect 2466 39686 2478 39738
rect 2478 39686 2492 39738
rect 2516 39686 2530 39738
rect 2530 39686 2542 39738
rect 2542 39686 2572 39738
rect 2596 39686 2606 39738
rect 2606 39686 2652 39738
rect 2356 39684 2412 39686
rect 2436 39684 2492 39686
rect 2516 39684 2572 39686
rect 2596 39684 2652 39686
rect 3016 39194 3072 39196
rect 3096 39194 3152 39196
rect 3176 39194 3232 39196
rect 3256 39194 3312 39196
rect 3016 39142 3062 39194
rect 3062 39142 3072 39194
rect 3096 39142 3126 39194
rect 3126 39142 3138 39194
rect 3138 39142 3152 39194
rect 3176 39142 3190 39194
rect 3190 39142 3202 39194
rect 3202 39142 3232 39194
rect 3256 39142 3266 39194
rect 3266 39142 3312 39194
rect 3016 39140 3072 39142
rect 3096 39140 3152 39142
rect 3176 39140 3232 39142
rect 3256 39140 3312 39142
rect 2356 38650 2412 38652
rect 2436 38650 2492 38652
rect 2516 38650 2572 38652
rect 2596 38650 2652 38652
rect 2356 38598 2402 38650
rect 2402 38598 2412 38650
rect 2436 38598 2466 38650
rect 2466 38598 2478 38650
rect 2478 38598 2492 38650
rect 2516 38598 2530 38650
rect 2530 38598 2542 38650
rect 2542 38598 2572 38650
rect 2596 38598 2606 38650
rect 2606 38598 2652 38650
rect 2356 38596 2412 38598
rect 2436 38596 2492 38598
rect 2516 38596 2572 38598
rect 2596 38596 2652 38598
rect 7356 45178 7412 45180
rect 7436 45178 7492 45180
rect 7516 45178 7572 45180
rect 7596 45178 7652 45180
rect 7356 45126 7402 45178
rect 7402 45126 7412 45178
rect 7436 45126 7466 45178
rect 7466 45126 7478 45178
rect 7478 45126 7492 45178
rect 7516 45126 7530 45178
rect 7530 45126 7542 45178
rect 7542 45126 7572 45178
rect 7596 45126 7606 45178
rect 7606 45126 7652 45178
rect 7356 45124 7412 45126
rect 7436 45124 7492 45126
rect 7516 45124 7572 45126
rect 7596 45124 7652 45126
rect 7356 44090 7412 44092
rect 7436 44090 7492 44092
rect 7516 44090 7572 44092
rect 7596 44090 7652 44092
rect 7356 44038 7402 44090
rect 7402 44038 7412 44090
rect 7436 44038 7466 44090
rect 7466 44038 7478 44090
rect 7478 44038 7492 44090
rect 7516 44038 7530 44090
rect 7530 44038 7542 44090
rect 7542 44038 7572 44090
rect 7596 44038 7606 44090
rect 7606 44038 7652 44090
rect 7356 44036 7412 44038
rect 7436 44036 7492 44038
rect 7516 44036 7572 44038
rect 7596 44036 7652 44038
rect 7356 43002 7412 43004
rect 7436 43002 7492 43004
rect 7516 43002 7572 43004
rect 7596 43002 7652 43004
rect 7356 42950 7402 43002
rect 7402 42950 7412 43002
rect 7436 42950 7466 43002
rect 7466 42950 7478 43002
rect 7478 42950 7492 43002
rect 7516 42950 7530 43002
rect 7530 42950 7542 43002
rect 7542 42950 7572 43002
rect 7596 42950 7606 43002
rect 7606 42950 7652 43002
rect 7356 42948 7412 42950
rect 7436 42948 7492 42950
rect 7516 42948 7572 42950
rect 7596 42948 7652 42950
rect 8016 47898 8072 47900
rect 8096 47898 8152 47900
rect 8176 47898 8232 47900
rect 8256 47898 8312 47900
rect 8016 47846 8062 47898
rect 8062 47846 8072 47898
rect 8096 47846 8126 47898
rect 8126 47846 8138 47898
rect 8138 47846 8152 47898
rect 8176 47846 8190 47898
rect 8190 47846 8202 47898
rect 8202 47846 8232 47898
rect 8256 47846 8266 47898
rect 8266 47846 8312 47898
rect 8016 47844 8072 47846
rect 8096 47844 8152 47846
rect 8176 47844 8232 47846
rect 8256 47844 8312 47846
rect 8390 47368 8446 47424
rect 8016 46810 8072 46812
rect 8096 46810 8152 46812
rect 8176 46810 8232 46812
rect 8256 46810 8312 46812
rect 8016 46758 8062 46810
rect 8062 46758 8072 46810
rect 8096 46758 8126 46810
rect 8126 46758 8138 46810
rect 8138 46758 8152 46810
rect 8176 46758 8190 46810
rect 8190 46758 8202 46810
rect 8202 46758 8232 46810
rect 8256 46758 8266 46810
rect 8266 46758 8312 46810
rect 8016 46756 8072 46758
rect 8096 46756 8152 46758
rect 8176 46756 8232 46758
rect 8256 46756 8312 46758
rect 8390 46008 8446 46064
rect 8016 45722 8072 45724
rect 8096 45722 8152 45724
rect 8176 45722 8232 45724
rect 8256 45722 8312 45724
rect 8016 45670 8062 45722
rect 8062 45670 8072 45722
rect 8096 45670 8126 45722
rect 8126 45670 8138 45722
rect 8138 45670 8152 45722
rect 8176 45670 8190 45722
rect 8190 45670 8202 45722
rect 8202 45670 8232 45722
rect 8256 45670 8266 45722
rect 8266 45670 8312 45722
rect 8016 45668 8072 45670
rect 8096 45668 8152 45670
rect 8176 45668 8232 45670
rect 8256 45668 8312 45670
rect 8390 44648 8446 44704
rect 8016 44634 8072 44636
rect 8096 44634 8152 44636
rect 8176 44634 8232 44636
rect 8256 44634 8312 44636
rect 8016 44582 8062 44634
rect 8062 44582 8072 44634
rect 8096 44582 8126 44634
rect 8126 44582 8138 44634
rect 8138 44582 8152 44634
rect 8176 44582 8190 44634
rect 8190 44582 8202 44634
rect 8202 44582 8232 44634
rect 8256 44582 8266 44634
rect 8266 44582 8312 44634
rect 8016 44580 8072 44582
rect 8096 44580 8152 44582
rect 8176 44580 8232 44582
rect 8256 44580 8312 44582
rect 8016 43546 8072 43548
rect 8096 43546 8152 43548
rect 8176 43546 8232 43548
rect 8256 43546 8312 43548
rect 8016 43494 8062 43546
rect 8062 43494 8072 43546
rect 8096 43494 8126 43546
rect 8126 43494 8138 43546
rect 8138 43494 8152 43546
rect 8176 43494 8190 43546
rect 8190 43494 8202 43546
rect 8202 43494 8232 43546
rect 8256 43494 8266 43546
rect 8266 43494 8312 43546
rect 8016 43492 8072 43494
rect 8096 43492 8152 43494
rect 8176 43492 8232 43494
rect 8256 43492 8312 43494
rect 8850 43288 8906 43344
rect 8016 42458 8072 42460
rect 8096 42458 8152 42460
rect 8176 42458 8232 42460
rect 8256 42458 8312 42460
rect 8016 42406 8062 42458
rect 8062 42406 8072 42458
rect 8096 42406 8126 42458
rect 8126 42406 8138 42458
rect 8138 42406 8152 42458
rect 8176 42406 8190 42458
rect 8190 42406 8202 42458
rect 8202 42406 8232 42458
rect 8256 42406 8266 42458
rect 8266 42406 8312 42458
rect 8016 42404 8072 42406
rect 8096 42404 8152 42406
rect 8176 42404 8232 42406
rect 8256 42404 8312 42406
rect 8390 41928 8446 41984
rect 7356 41914 7412 41916
rect 7436 41914 7492 41916
rect 7516 41914 7572 41916
rect 7596 41914 7652 41916
rect 7356 41862 7402 41914
rect 7402 41862 7412 41914
rect 7436 41862 7466 41914
rect 7466 41862 7478 41914
rect 7478 41862 7492 41914
rect 7516 41862 7530 41914
rect 7530 41862 7542 41914
rect 7542 41862 7572 41914
rect 7596 41862 7606 41914
rect 7606 41862 7652 41914
rect 7356 41860 7412 41862
rect 7436 41860 7492 41862
rect 7516 41860 7572 41862
rect 7596 41860 7652 41862
rect 7356 40826 7412 40828
rect 7436 40826 7492 40828
rect 7516 40826 7572 40828
rect 7596 40826 7652 40828
rect 7356 40774 7402 40826
rect 7402 40774 7412 40826
rect 7436 40774 7466 40826
rect 7466 40774 7478 40826
rect 7478 40774 7492 40826
rect 7516 40774 7530 40826
rect 7530 40774 7542 40826
rect 7542 40774 7572 40826
rect 7596 40774 7606 40826
rect 7606 40774 7652 40826
rect 7356 40772 7412 40774
rect 7436 40772 7492 40774
rect 7516 40772 7572 40774
rect 7596 40772 7652 40774
rect 3016 38106 3072 38108
rect 3096 38106 3152 38108
rect 3176 38106 3232 38108
rect 3256 38106 3312 38108
rect 3016 38054 3062 38106
rect 3062 38054 3072 38106
rect 3096 38054 3126 38106
rect 3126 38054 3138 38106
rect 3138 38054 3152 38106
rect 3176 38054 3190 38106
rect 3190 38054 3202 38106
rect 3202 38054 3232 38106
rect 3256 38054 3266 38106
rect 3266 38054 3312 38106
rect 3016 38052 3072 38054
rect 3096 38052 3152 38054
rect 3176 38052 3232 38054
rect 3256 38052 3312 38054
rect 2356 37562 2412 37564
rect 2436 37562 2492 37564
rect 2516 37562 2572 37564
rect 2596 37562 2652 37564
rect 2356 37510 2402 37562
rect 2402 37510 2412 37562
rect 2436 37510 2466 37562
rect 2466 37510 2478 37562
rect 2478 37510 2492 37562
rect 2516 37510 2530 37562
rect 2530 37510 2542 37562
rect 2542 37510 2572 37562
rect 2596 37510 2606 37562
rect 2606 37510 2652 37562
rect 2356 37508 2412 37510
rect 2436 37508 2492 37510
rect 2516 37508 2572 37510
rect 2596 37508 2652 37510
rect 3016 37018 3072 37020
rect 3096 37018 3152 37020
rect 3176 37018 3232 37020
rect 3256 37018 3312 37020
rect 3016 36966 3062 37018
rect 3062 36966 3072 37018
rect 3096 36966 3126 37018
rect 3126 36966 3138 37018
rect 3138 36966 3152 37018
rect 3176 36966 3190 37018
rect 3190 36966 3202 37018
rect 3202 36966 3232 37018
rect 3256 36966 3266 37018
rect 3266 36966 3312 37018
rect 3016 36964 3072 36966
rect 3096 36964 3152 36966
rect 3176 36964 3232 36966
rect 3256 36964 3312 36966
rect 2356 36474 2412 36476
rect 2436 36474 2492 36476
rect 2516 36474 2572 36476
rect 2596 36474 2652 36476
rect 2356 36422 2402 36474
rect 2402 36422 2412 36474
rect 2436 36422 2466 36474
rect 2466 36422 2478 36474
rect 2478 36422 2492 36474
rect 2516 36422 2530 36474
rect 2530 36422 2542 36474
rect 2542 36422 2572 36474
rect 2596 36422 2606 36474
rect 2606 36422 2652 36474
rect 2356 36420 2412 36422
rect 2436 36420 2492 36422
rect 2516 36420 2572 36422
rect 2596 36420 2652 36422
rect 3016 35930 3072 35932
rect 3096 35930 3152 35932
rect 3176 35930 3232 35932
rect 3256 35930 3312 35932
rect 3016 35878 3062 35930
rect 3062 35878 3072 35930
rect 3096 35878 3126 35930
rect 3126 35878 3138 35930
rect 3138 35878 3152 35930
rect 3176 35878 3190 35930
rect 3190 35878 3202 35930
rect 3202 35878 3232 35930
rect 3256 35878 3266 35930
rect 3266 35878 3312 35930
rect 3016 35876 3072 35878
rect 3096 35876 3152 35878
rect 3176 35876 3232 35878
rect 3256 35876 3312 35878
rect 2356 35386 2412 35388
rect 2436 35386 2492 35388
rect 2516 35386 2572 35388
rect 2596 35386 2652 35388
rect 2356 35334 2402 35386
rect 2402 35334 2412 35386
rect 2436 35334 2466 35386
rect 2466 35334 2478 35386
rect 2478 35334 2492 35386
rect 2516 35334 2530 35386
rect 2530 35334 2542 35386
rect 2542 35334 2572 35386
rect 2596 35334 2606 35386
rect 2606 35334 2652 35386
rect 2356 35332 2412 35334
rect 2436 35332 2492 35334
rect 2516 35332 2572 35334
rect 2596 35332 2652 35334
rect 3016 34842 3072 34844
rect 3096 34842 3152 34844
rect 3176 34842 3232 34844
rect 3256 34842 3312 34844
rect 3016 34790 3062 34842
rect 3062 34790 3072 34842
rect 3096 34790 3126 34842
rect 3126 34790 3138 34842
rect 3138 34790 3152 34842
rect 3176 34790 3190 34842
rect 3190 34790 3202 34842
rect 3202 34790 3232 34842
rect 3256 34790 3266 34842
rect 3266 34790 3312 34842
rect 3016 34788 3072 34790
rect 3096 34788 3152 34790
rect 3176 34788 3232 34790
rect 3256 34788 3312 34790
rect 2356 34298 2412 34300
rect 2436 34298 2492 34300
rect 2516 34298 2572 34300
rect 2596 34298 2652 34300
rect 2356 34246 2402 34298
rect 2402 34246 2412 34298
rect 2436 34246 2466 34298
rect 2466 34246 2478 34298
rect 2478 34246 2492 34298
rect 2516 34246 2530 34298
rect 2530 34246 2542 34298
rect 2542 34246 2572 34298
rect 2596 34246 2606 34298
rect 2606 34246 2652 34298
rect 2356 34244 2412 34246
rect 2436 34244 2492 34246
rect 2516 34244 2572 34246
rect 2596 34244 2652 34246
rect 3016 33754 3072 33756
rect 3096 33754 3152 33756
rect 3176 33754 3232 33756
rect 3256 33754 3312 33756
rect 3016 33702 3062 33754
rect 3062 33702 3072 33754
rect 3096 33702 3126 33754
rect 3126 33702 3138 33754
rect 3138 33702 3152 33754
rect 3176 33702 3190 33754
rect 3190 33702 3202 33754
rect 3202 33702 3232 33754
rect 3256 33702 3266 33754
rect 3266 33702 3312 33754
rect 3016 33700 3072 33702
rect 3096 33700 3152 33702
rect 3176 33700 3232 33702
rect 3256 33700 3312 33702
rect 2356 33210 2412 33212
rect 2436 33210 2492 33212
rect 2516 33210 2572 33212
rect 2596 33210 2652 33212
rect 2356 33158 2402 33210
rect 2402 33158 2412 33210
rect 2436 33158 2466 33210
rect 2466 33158 2478 33210
rect 2478 33158 2492 33210
rect 2516 33158 2530 33210
rect 2530 33158 2542 33210
rect 2542 33158 2572 33210
rect 2596 33158 2606 33210
rect 2606 33158 2652 33210
rect 2356 33156 2412 33158
rect 2436 33156 2492 33158
rect 2516 33156 2572 33158
rect 2596 33156 2652 33158
rect 3016 32666 3072 32668
rect 3096 32666 3152 32668
rect 3176 32666 3232 32668
rect 3256 32666 3312 32668
rect 3016 32614 3062 32666
rect 3062 32614 3072 32666
rect 3096 32614 3126 32666
rect 3126 32614 3138 32666
rect 3138 32614 3152 32666
rect 3176 32614 3190 32666
rect 3190 32614 3202 32666
rect 3202 32614 3232 32666
rect 3256 32614 3266 32666
rect 3266 32614 3312 32666
rect 3016 32612 3072 32614
rect 3096 32612 3152 32614
rect 3176 32612 3232 32614
rect 3256 32612 3312 32614
rect 2356 32122 2412 32124
rect 2436 32122 2492 32124
rect 2516 32122 2572 32124
rect 2596 32122 2652 32124
rect 2356 32070 2402 32122
rect 2402 32070 2412 32122
rect 2436 32070 2466 32122
rect 2466 32070 2478 32122
rect 2478 32070 2492 32122
rect 2516 32070 2530 32122
rect 2530 32070 2542 32122
rect 2542 32070 2572 32122
rect 2596 32070 2606 32122
rect 2606 32070 2652 32122
rect 2356 32068 2412 32070
rect 2436 32068 2492 32070
rect 2516 32068 2572 32070
rect 2596 32068 2652 32070
rect 3016 31578 3072 31580
rect 3096 31578 3152 31580
rect 3176 31578 3232 31580
rect 3256 31578 3312 31580
rect 3016 31526 3062 31578
rect 3062 31526 3072 31578
rect 3096 31526 3126 31578
rect 3126 31526 3138 31578
rect 3138 31526 3152 31578
rect 3176 31526 3190 31578
rect 3190 31526 3202 31578
rect 3202 31526 3232 31578
rect 3256 31526 3266 31578
rect 3266 31526 3312 31578
rect 3016 31524 3072 31526
rect 3096 31524 3152 31526
rect 3176 31524 3232 31526
rect 3256 31524 3312 31526
rect 2356 31034 2412 31036
rect 2436 31034 2492 31036
rect 2516 31034 2572 31036
rect 2596 31034 2652 31036
rect 2356 30982 2402 31034
rect 2402 30982 2412 31034
rect 2436 30982 2466 31034
rect 2466 30982 2478 31034
rect 2478 30982 2492 31034
rect 2516 30982 2530 31034
rect 2530 30982 2542 31034
rect 2542 30982 2572 31034
rect 2596 30982 2606 31034
rect 2606 30982 2652 31034
rect 2356 30980 2412 30982
rect 2436 30980 2492 30982
rect 2516 30980 2572 30982
rect 2596 30980 2652 30982
rect 3016 30490 3072 30492
rect 3096 30490 3152 30492
rect 3176 30490 3232 30492
rect 3256 30490 3312 30492
rect 3016 30438 3062 30490
rect 3062 30438 3072 30490
rect 3096 30438 3126 30490
rect 3126 30438 3138 30490
rect 3138 30438 3152 30490
rect 3176 30438 3190 30490
rect 3190 30438 3202 30490
rect 3202 30438 3232 30490
rect 3256 30438 3266 30490
rect 3266 30438 3312 30490
rect 3016 30436 3072 30438
rect 3096 30436 3152 30438
rect 3176 30436 3232 30438
rect 3256 30436 3312 30438
rect 2356 29946 2412 29948
rect 2436 29946 2492 29948
rect 2516 29946 2572 29948
rect 2596 29946 2652 29948
rect 2356 29894 2402 29946
rect 2402 29894 2412 29946
rect 2436 29894 2466 29946
rect 2466 29894 2478 29946
rect 2478 29894 2492 29946
rect 2516 29894 2530 29946
rect 2530 29894 2542 29946
rect 2542 29894 2572 29946
rect 2596 29894 2606 29946
rect 2606 29894 2652 29946
rect 2356 29892 2412 29894
rect 2436 29892 2492 29894
rect 2516 29892 2572 29894
rect 2596 29892 2652 29894
rect 3016 29402 3072 29404
rect 3096 29402 3152 29404
rect 3176 29402 3232 29404
rect 3256 29402 3312 29404
rect 3016 29350 3062 29402
rect 3062 29350 3072 29402
rect 3096 29350 3126 29402
rect 3126 29350 3138 29402
rect 3138 29350 3152 29402
rect 3176 29350 3190 29402
rect 3190 29350 3202 29402
rect 3202 29350 3232 29402
rect 3256 29350 3266 29402
rect 3266 29350 3312 29402
rect 3016 29348 3072 29350
rect 3096 29348 3152 29350
rect 3176 29348 3232 29350
rect 3256 29348 3312 29350
rect 2356 28858 2412 28860
rect 2436 28858 2492 28860
rect 2516 28858 2572 28860
rect 2596 28858 2652 28860
rect 2356 28806 2402 28858
rect 2402 28806 2412 28858
rect 2436 28806 2466 28858
rect 2466 28806 2478 28858
rect 2478 28806 2492 28858
rect 2516 28806 2530 28858
rect 2530 28806 2542 28858
rect 2542 28806 2572 28858
rect 2596 28806 2606 28858
rect 2606 28806 2652 28858
rect 2356 28804 2412 28806
rect 2436 28804 2492 28806
rect 2516 28804 2572 28806
rect 2596 28804 2652 28806
rect 3016 28314 3072 28316
rect 3096 28314 3152 28316
rect 3176 28314 3232 28316
rect 3256 28314 3312 28316
rect 3016 28262 3062 28314
rect 3062 28262 3072 28314
rect 3096 28262 3126 28314
rect 3126 28262 3138 28314
rect 3138 28262 3152 28314
rect 3176 28262 3190 28314
rect 3190 28262 3202 28314
rect 3202 28262 3232 28314
rect 3256 28262 3266 28314
rect 3266 28262 3312 28314
rect 3016 28260 3072 28262
rect 3096 28260 3152 28262
rect 3176 28260 3232 28262
rect 3256 28260 3312 28262
rect 2356 27770 2412 27772
rect 2436 27770 2492 27772
rect 2516 27770 2572 27772
rect 2596 27770 2652 27772
rect 2356 27718 2402 27770
rect 2402 27718 2412 27770
rect 2436 27718 2466 27770
rect 2466 27718 2478 27770
rect 2478 27718 2492 27770
rect 2516 27718 2530 27770
rect 2530 27718 2542 27770
rect 2542 27718 2572 27770
rect 2596 27718 2606 27770
rect 2606 27718 2652 27770
rect 2356 27716 2412 27718
rect 2436 27716 2492 27718
rect 2516 27716 2572 27718
rect 2596 27716 2652 27718
rect 3016 27226 3072 27228
rect 3096 27226 3152 27228
rect 3176 27226 3232 27228
rect 3256 27226 3312 27228
rect 3016 27174 3062 27226
rect 3062 27174 3072 27226
rect 3096 27174 3126 27226
rect 3126 27174 3138 27226
rect 3138 27174 3152 27226
rect 3176 27174 3190 27226
rect 3190 27174 3202 27226
rect 3202 27174 3232 27226
rect 3256 27174 3266 27226
rect 3266 27174 3312 27226
rect 3016 27172 3072 27174
rect 3096 27172 3152 27174
rect 3176 27172 3232 27174
rect 3256 27172 3312 27174
rect 2356 26682 2412 26684
rect 2436 26682 2492 26684
rect 2516 26682 2572 26684
rect 2596 26682 2652 26684
rect 2356 26630 2402 26682
rect 2402 26630 2412 26682
rect 2436 26630 2466 26682
rect 2466 26630 2478 26682
rect 2478 26630 2492 26682
rect 2516 26630 2530 26682
rect 2530 26630 2542 26682
rect 2542 26630 2572 26682
rect 2596 26630 2606 26682
rect 2606 26630 2652 26682
rect 2356 26628 2412 26630
rect 2436 26628 2492 26630
rect 2516 26628 2572 26630
rect 2596 26628 2652 26630
rect 3016 26138 3072 26140
rect 3096 26138 3152 26140
rect 3176 26138 3232 26140
rect 3256 26138 3312 26140
rect 3016 26086 3062 26138
rect 3062 26086 3072 26138
rect 3096 26086 3126 26138
rect 3126 26086 3138 26138
rect 3138 26086 3152 26138
rect 3176 26086 3190 26138
rect 3190 26086 3202 26138
rect 3202 26086 3232 26138
rect 3256 26086 3266 26138
rect 3266 26086 3312 26138
rect 3016 26084 3072 26086
rect 3096 26084 3152 26086
rect 3176 26084 3232 26086
rect 3256 26084 3312 26086
rect 2356 25594 2412 25596
rect 2436 25594 2492 25596
rect 2516 25594 2572 25596
rect 2596 25594 2652 25596
rect 2356 25542 2402 25594
rect 2402 25542 2412 25594
rect 2436 25542 2466 25594
rect 2466 25542 2478 25594
rect 2478 25542 2492 25594
rect 2516 25542 2530 25594
rect 2530 25542 2542 25594
rect 2542 25542 2572 25594
rect 2596 25542 2606 25594
rect 2606 25542 2652 25594
rect 2356 25540 2412 25542
rect 2436 25540 2492 25542
rect 2516 25540 2572 25542
rect 2596 25540 2652 25542
rect 3016 25050 3072 25052
rect 3096 25050 3152 25052
rect 3176 25050 3232 25052
rect 3256 25050 3312 25052
rect 3016 24998 3062 25050
rect 3062 24998 3072 25050
rect 3096 24998 3126 25050
rect 3126 24998 3138 25050
rect 3138 24998 3152 25050
rect 3176 24998 3190 25050
rect 3190 24998 3202 25050
rect 3202 24998 3232 25050
rect 3256 24998 3266 25050
rect 3266 24998 3312 25050
rect 3016 24996 3072 24998
rect 3096 24996 3152 24998
rect 3176 24996 3232 24998
rect 3256 24996 3312 24998
rect 2356 24506 2412 24508
rect 2436 24506 2492 24508
rect 2516 24506 2572 24508
rect 2596 24506 2652 24508
rect 2356 24454 2402 24506
rect 2402 24454 2412 24506
rect 2436 24454 2466 24506
rect 2466 24454 2478 24506
rect 2478 24454 2492 24506
rect 2516 24454 2530 24506
rect 2530 24454 2542 24506
rect 2542 24454 2572 24506
rect 2596 24454 2606 24506
rect 2606 24454 2652 24506
rect 2356 24452 2412 24454
rect 2436 24452 2492 24454
rect 2516 24452 2572 24454
rect 2596 24452 2652 24454
rect 7356 39738 7412 39740
rect 7436 39738 7492 39740
rect 7516 39738 7572 39740
rect 7596 39738 7652 39740
rect 7356 39686 7402 39738
rect 7402 39686 7412 39738
rect 7436 39686 7466 39738
rect 7466 39686 7478 39738
rect 7478 39686 7492 39738
rect 7516 39686 7530 39738
rect 7530 39686 7542 39738
rect 7542 39686 7572 39738
rect 7596 39686 7606 39738
rect 7606 39686 7652 39738
rect 7356 39684 7412 39686
rect 7436 39684 7492 39686
rect 7516 39684 7572 39686
rect 7596 39684 7652 39686
rect 7356 38650 7412 38652
rect 7436 38650 7492 38652
rect 7516 38650 7572 38652
rect 7596 38650 7652 38652
rect 7356 38598 7402 38650
rect 7402 38598 7412 38650
rect 7436 38598 7466 38650
rect 7466 38598 7478 38650
rect 7478 38598 7492 38650
rect 7516 38598 7530 38650
rect 7530 38598 7542 38650
rect 7542 38598 7572 38650
rect 7596 38598 7606 38650
rect 7606 38598 7652 38650
rect 7356 38596 7412 38598
rect 7436 38596 7492 38598
rect 7516 38596 7572 38598
rect 7596 38596 7652 38598
rect 7356 37562 7412 37564
rect 7436 37562 7492 37564
rect 7516 37562 7572 37564
rect 7596 37562 7652 37564
rect 7356 37510 7402 37562
rect 7402 37510 7412 37562
rect 7436 37510 7466 37562
rect 7466 37510 7478 37562
rect 7478 37510 7492 37562
rect 7516 37510 7530 37562
rect 7530 37510 7542 37562
rect 7542 37510 7572 37562
rect 7596 37510 7606 37562
rect 7606 37510 7652 37562
rect 7356 37508 7412 37510
rect 7436 37508 7492 37510
rect 7516 37508 7572 37510
rect 7596 37508 7652 37510
rect 7356 36474 7412 36476
rect 7436 36474 7492 36476
rect 7516 36474 7572 36476
rect 7596 36474 7652 36476
rect 7356 36422 7402 36474
rect 7402 36422 7412 36474
rect 7436 36422 7466 36474
rect 7466 36422 7478 36474
rect 7478 36422 7492 36474
rect 7516 36422 7530 36474
rect 7530 36422 7542 36474
rect 7542 36422 7572 36474
rect 7596 36422 7606 36474
rect 7606 36422 7652 36474
rect 7356 36420 7412 36422
rect 7436 36420 7492 36422
rect 7516 36420 7572 36422
rect 7596 36420 7652 36422
rect 3016 23962 3072 23964
rect 3096 23962 3152 23964
rect 3176 23962 3232 23964
rect 3256 23962 3312 23964
rect 3016 23910 3062 23962
rect 3062 23910 3072 23962
rect 3096 23910 3126 23962
rect 3126 23910 3138 23962
rect 3138 23910 3152 23962
rect 3176 23910 3190 23962
rect 3190 23910 3202 23962
rect 3202 23910 3232 23962
rect 3256 23910 3266 23962
rect 3266 23910 3312 23962
rect 3016 23908 3072 23910
rect 3096 23908 3152 23910
rect 3176 23908 3232 23910
rect 3256 23908 3312 23910
rect 2356 23418 2412 23420
rect 2436 23418 2492 23420
rect 2516 23418 2572 23420
rect 2596 23418 2652 23420
rect 2356 23366 2402 23418
rect 2402 23366 2412 23418
rect 2436 23366 2466 23418
rect 2466 23366 2478 23418
rect 2478 23366 2492 23418
rect 2516 23366 2530 23418
rect 2530 23366 2542 23418
rect 2542 23366 2572 23418
rect 2596 23366 2606 23418
rect 2606 23366 2652 23418
rect 2356 23364 2412 23366
rect 2436 23364 2492 23366
rect 2516 23364 2572 23366
rect 2596 23364 2652 23366
rect 3016 22874 3072 22876
rect 3096 22874 3152 22876
rect 3176 22874 3232 22876
rect 3256 22874 3312 22876
rect 3016 22822 3062 22874
rect 3062 22822 3072 22874
rect 3096 22822 3126 22874
rect 3126 22822 3138 22874
rect 3138 22822 3152 22874
rect 3176 22822 3190 22874
rect 3190 22822 3202 22874
rect 3202 22822 3232 22874
rect 3256 22822 3266 22874
rect 3266 22822 3312 22874
rect 3016 22820 3072 22822
rect 3096 22820 3152 22822
rect 3176 22820 3232 22822
rect 3256 22820 3312 22822
rect 2356 22330 2412 22332
rect 2436 22330 2492 22332
rect 2516 22330 2572 22332
rect 2596 22330 2652 22332
rect 2356 22278 2402 22330
rect 2402 22278 2412 22330
rect 2436 22278 2466 22330
rect 2466 22278 2478 22330
rect 2478 22278 2492 22330
rect 2516 22278 2530 22330
rect 2530 22278 2542 22330
rect 2542 22278 2572 22330
rect 2596 22278 2606 22330
rect 2606 22278 2652 22330
rect 2356 22276 2412 22278
rect 2436 22276 2492 22278
rect 2516 22276 2572 22278
rect 2596 22276 2652 22278
rect 3016 21786 3072 21788
rect 3096 21786 3152 21788
rect 3176 21786 3232 21788
rect 3256 21786 3312 21788
rect 3016 21734 3062 21786
rect 3062 21734 3072 21786
rect 3096 21734 3126 21786
rect 3126 21734 3138 21786
rect 3138 21734 3152 21786
rect 3176 21734 3190 21786
rect 3190 21734 3202 21786
rect 3202 21734 3232 21786
rect 3256 21734 3266 21786
rect 3266 21734 3312 21786
rect 3016 21732 3072 21734
rect 3096 21732 3152 21734
rect 3176 21732 3232 21734
rect 3256 21732 3312 21734
rect 2356 21242 2412 21244
rect 2436 21242 2492 21244
rect 2516 21242 2572 21244
rect 2596 21242 2652 21244
rect 2356 21190 2402 21242
rect 2402 21190 2412 21242
rect 2436 21190 2466 21242
rect 2466 21190 2478 21242
rect 2478 21190 2492 21242
rect 2516 21190 2530 21242
rect 2530 21190 2542 21242
rect 2542 21190 2572 21242
rect 2596 21190 2606 21242
rect 2606 21190 2652 21242
rect 2356 21188 2412 21190
rect 2436 21188 2492 21190
rect 2516 21188 2572 21190
rect 2596 21188 2652 21190
rect 3016 20698 3072 20700
rect 3096 20698 3152 20700
rect 3176 20698 3232 20700
rect 3256 20698 3312 20700
rect 3016 20646 3062 20698
rect 3062 20646 3072 20698
rect 3096 20646 3126 20698
rect 3126 20646 3138 20698
rect 3138 20646 3152 20698
rect 3176 20646 3190 20698
rect 3190 20646 3202 20698
rect 3202 20646 3232 20698
rect 3256 20646 3266 20698
rect 3266 20646 3312 20698
rect 3016 20644 3072 20646
rect 3096 20644 3152 20646
rect 3176 20644 3232 20646
rect 3256 20644 3312 20646
rect 2356 20154 2412 20156
rect 2436 20154 2492 20156
rect 2516 20154 2572 20156
rect 2596 20154 2652 20156
rect 2356 20102 2402 20154
rect 2402 20102 2412 20154
rect 2436 20102 2466 20154
rect 2466 20102 2478 20154
rect 2478 20102 2492 20154
rect 2516 20102 2530 20154
rect 2530 20102 2542 20154
rect 2542 20102 2572 20154
rect 2596 20102 2606 20154
rect 2606 20102 2652 20154
rect 2356 20100 2412 20102
rect 2436 20100 2492 20102
rect 2516 20100 2572 20102
rect 2596 20100 2652 20102
rect 3016 19610 3072 19612
rect 3096 19610 3152 19612
rect 3176 19610 3232 19612
rect 3256 19610 3312 19612
rect 3016 19558 3062 19610
rect 3062 19558 3072 19610
rect 3096 19558 3126 19610
rect 3126 19558 3138 19610
rect 3138 19558 3152 19610
rect 3176 19558 3190 19610
rect 3190 19558 3202 19610
rect 3202 19558 3232 19610
rect 3256 19558 3266 19610
rect 3266 19558 3312 19610
rect 3016 19556 3072 19558
rect 3096 19556 3152 19558
rect 3176 19556 3232 19558
rect 3256 19556 3312 19558
rect 2356 19066 2412 19068
rect 2436 19066 2492 19068
rect 2516 19066 2572 19068
rect 2596 19066 2652 19068
rect 2356 19014 2402 19066
rect 2402 19014 2412 19066
rect 2436 19014 2466 19066
rect 2466 19014 2478 19066
rect 2478 19014 2492 19066
rect 2516 19014 2530 19066
rect 2530 19014 2542 19066
rect 2542 19014 2572 19066
rect 2596 19014 2606 19066
rect 2606 19014 2652 19066
rect 2356 19012 2412 19014
rect 2436 19012 2492 19014
rect 2516 19012 2572 19014
rect 2596 19012 2652 19014
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 3176 18522 3232 18524
rect 3256 18522 3312 18524
rect 3016 18470 3062 18522
rect 3062 18470 3072 18522
rect 3096 18470 3126 18522
rect 3126 18470 3138 18522
rect 3138 18470 3152 18522
rect 3176 18470 3190 18522
rect 3190 18470 3202 18522
rect 3202 18470 3232 18522
rect 3256 18470 3266 18522
rect 3266 18470 3312 18522
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 3176 18468 3232 18470
rect 3256 18468 3312 18470
rect 2356 17978 2412 17980
rect 2436 17978 2492 17980
rect 2516 17978 2572 17980
rect 2596 17978 2652 17980
rect 2356 17926 2402 17978
rect 2402 17926 2412 17978
rect 2436 17926 2466 17978
rect 2466 17926 2478 17978
rect 2478 17926 2492 17978
rect 2516 17926 2530 17978
rect 2530 17926 2542 17978
rect 2542 17926 2572 17978
rect 2596 17926 2606 17978
rect 2606 17926 2652 17978
rect 2356 17924 2412 17926
rect 2436 17924 2492 17926
rect 2516 17924 2572 17926
rect 2596 17924 2652 17926
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 3176 17434 3232 17436
rect 3256 17434 3312 17436
rect 3016 17382 3062 17434
rect 3062 17382 3072 17434
rect 3096 17382 3126 17434
rect 3126 17382 3138 17434
rect 3138 17382 3152 17434
rect 3176 17382 3190 17434
rect 3190 17382 3202 17434
rect 3202 17382 3232 17434
rect 3256 17382 3266 17434
rect 3266 17382 3312 17434
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 3176 17380 3232 17382
rect 3256 17380 3312 17382
rect 2356 16890 2412 16892
rect 2436 16890 2492 16892
rect 2516 16890 2572 16892
rect 2596 16890 2652 16892
rect 2356 16838 2402 16890
rect 2402 16838 2412 16890
rect 2436 16838 2466 16890
rect 2466 16838 2478 16890
rect 2478 16838 2492 16890
rect 2516 16838 2530 16890
rect 2530 16838 2542 16890
rect 2542 16838 2572 16890
rect 2596 16838 2606 16890
rect 2606 16838 2652 16890
rect 2356 16836 2412 16838
rect 2436 16836 2492 16838
rect 2516 16836 2572 16838
rect 2596 16836 2652 16838
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 3176 16346 3232 16348
rect 3256 16346 3312 16348
rect 3016 16294 3062 16346
rect 3062 16294 3072 16346
rect 3096 16294 3126 16346
rect 3126 16294 3138 16346
rect 3138 16294 3152 16346
rect 3176 16294 3190 16346
rect 3190 16294 3202 16346
rect 3202 16294 3232 16346
rect 3256 16294 3266 16346
rect 3266 16294 3312 16346
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 3176 16292 3232 16294
rect 3256 16292 3312 16294
rect 2356 15802 2412 15804
rect 2436 15802 2492 15804
rect 2516 15802 2572 15804
rect 2596 15802 2652 15804
rect 2356 15750 2402 15802
rect 2402 15750 2412 15802
rect 2436 15750 2466 15802
rect 2466 15750 2478 15802
rect 2478 15750 2492 15802
rect 2516 15750 2530 15802
rect 2530 15750 2542 15802
rect 2542 15750 2572 15802
rect 2596 15750 2606 15802
rect 2606 15750 2652 15802
rect 2356 15748 2412 15750
rect 2436 15748 2492 15750
rect 2516 15748 2572 15750
rect 2596 15748 2652 15750
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 3176 15258 3232 15260
rect 3256 15258 3312 15260
rect 3016 15206 3062 15258
rect 3062 15206 3072 15258
rect 3096 15206 3126 15258
rect 3126 15206 3138 15258
rect 3138 15206 3152 15258
rect 3176 15206 3190 15258
rect 3190 15206 3202 15258
rect 3202 15206 3232 15258
rect 3256 15206 3266 15258
rect 3266 15206 3312 15258
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 3176 15204 3232 15206
rect 3256 15204 3312 15206
rect 2356 14714 2412 14716
rect 2436 14714 2492 14716
rect 2516 14714 2572 14716
rect 2596 14714 2652 14716
rect 2356 14662 2402 14714
rect 2402 14662 2412 14714
rect 2436 14662 2466 14714
rect 2466 14662 2478 14714
rect 2478 14662 2492 14714
rect 2516 14662 2530 14714
rect 2530 14662 2542 14714
rect 2542 14662 2572 14714
rect 2596 14662 2606 14714
rect 2606 14662 2652 14714
rect 2356 14660 2412 14662
rect 2436 14660 2492 14662
rect 2516 14660 2572 14662
rect 2596 14660 2652 14662
rect 6734 16088 6790 16144
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 3176 14170 3232 14172
rect 3256 14170 3312 14172
rect 3016 14118 3062 14170
rect 3062 14118 3072 14170
rect 3096 14118 3126 14170
rect 3126 14118 3138 14170
rect 3138 14118 3152 14170
rect 3176 14118 3190 14170
rect 3190 14118 3202 14170
rect 3202 14118 3232 14170
rect 3256 14118 3266 14170
rect 3266 14118 3312 14170
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 3176 14116 3232 14118
rect 3256 14116 3312 14118
rect 2356 13626 2412 13628
rect 2436 13626 2492 13628
rect 2516 13626 2572 13628
rect 2596 13626 2652 13628
rect 2356 13574 2402 13626
rect 2402 13574 2412 13626
rect 2436 13574 2466 13626
rect 2466 13574 2478 13626
rect 2478 13574 2492 13626
rect 2516 13574 2530 13626
rect 2530 13574 2542 13626
rect 2542 13574 2572 13626
rect 2596 13574 2606 13626
rect 2606 13574 2652 13626
rect 2356 13572 2412 13574
rect 2436 13572 2492 13574
rect 2516 13572 2572 13574
rect 2596 13572 2652 13574
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 3176 13082 3232 13084
rect 3256 13082 3312 13084
rect 3016 13030 3062 13082
rect 3062 13030 3072 13082
rect 3096 13030 3126 13082
rect 3126 13030 3138 13082
rect 3138 13030 3152 13082
rect 3176 13030 3190 13082
rect 3190 13030 3202 13082
rect 3202 13030 3232 13082
rect 3256 13030 3266 13082
rect 3266 13030 3312 13082
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 3176 13028 3232 13030
rect 3256 13028 3312 13030
rect 7356 35386 7412 35388
rect 7436 35386 7492 35388
rect 7516 35386 7572 35388
rect 7596 35386 7652 35388
rect 7356 35334 7402 35386
rect 7402 35334 7412 35386
rect 7436 35334 7466 35386
rect 7466 35334 7478 35386
rect 7478 35334 7492 35386
rect 7516 35334 7530 35386
rect 7530 35334 7542 35386
rect 7542 35334 7572 35386
rect 7596 35334 7606 35386
rect 7606 35334 7652 35386
rect 7356 35332 7412 35334
rect 7436 35332 7492 35334
rect 7516 35332 7572 35334
rect 7596 35332 7652 35334
rect 7356 34298 7412 34300
rect 7436 34298 7492 34300
rect 7516 34298 7572 34300
rect 7596 34298 7652 34300
rect 7356 34246 7402 34298
rect 7402 34246 7412 34298
rect 7436 34246 7466 34298
rect 7466 34246 7478 34298
rect 7478 34246 7492 34298
rect 7516 34246 7530 34298
rect 7530 34246 7542 34298
rect 7542 34246 7572 34298
rect 7596 34246 7606 34298
rect 7606 34246 7652 34298
rect 7356 34244 7412 34246
rect 7436 34244 7492 34246
rect 7516 34244 7572 34246
rect 7596 34244 7652 34246
rect 7746 33496 7802 33552
rect 7356 33210 7412 33212
rect 7436 33210 7492 33212
rect 7516 33210 7572 33212
rect 7596 33210 7652 33212
rect 7356 33158 7402 33210
rect 7402 33158 7412 33210
rect 7436 33158 7466 33210
rect 7466 33158 7478 33210
rect 7478 33158 7492 33210
rect 7516 33158 7530 33210
rect 7530 33158 7542 33210
rect 7542 33158 7572 33210
rect 7596 33158 7606 33210
rect 7606 33158 7652 33210
rect 7356 33156 7412 33158
rect 7436 33156 7492 33158
rect 7516 33156 7572 33158
rect 7596 33156 7652 33158
rect 7356 32122 7412 32124
rect 7436 32122 7492 32124
rect 7516 32122 7572 32124
rect 7596 32122 7652 32124
rect 7356 32070 7402 32122
rect 7402 32070 7412 32122
rect 7436 32070 7466 32122
rect 7466 32070 7478 32122
rect 7478 32070 7492 32122
rect 7516 32070 7530 32122
rect 7530 32070 7542 32122
rect 7542 32070 7572 32122
rect 7596 32070 7606 32122
rect 7606 32070 7652 32122
rect 7356 32068 7412 32070
rect 7436 32068 7492 32070
rect 7516 32068 7572 32070
rect 7596 32068 7652 32070
rect 7356 31034 7412 31036
rect 7436 31034 7492 31036
rect 7516 31034 7572 31036
rect 7596 31034 7652 31036
rect 7356 30982 7402 31034
rect 7402 30982 7412 31034
rect 7436 30982 7466 31034
rect 7466 30982 7478 31034
rect 7478 30982 7492 31034
rect 7516 30982 7530 31034
rect 7530 30982 7542 31034
rect 7542 30982 7572 31034
rect 7596 30982 7606 31034
rect 7606 30982 7652 31034
rect 7356 30980 7412 30982
rect 7436 30980 7492 30982
rect 7516 30980 7572 30982
rect 7596 30980 7652 30982
rect 7356 29946 7412 29948
rect 7436 29946 7492 29948
rect 7516 29946 7572 29948
rect 7596 29946 7652 29948
rect 7356 29894 7402 29946
rect 7402 29894 7412 29946
rect 7436 29894 7466 29946
rect 7466 29894 7478 29946
rect 7478 29894 7492 29946
rect 7516 29894 7530 29946
rect 7530 29894 7542 29946
rect 7542 29894 7572 29946
rect 7596 29894 7606 29946
rect 7606 29894 7652 29946
rect 7356 29892 7412 29894
rect 7436 29892 7492 29894
rect 7516 29892 7572 29894
rect 7596 29892 7652 29894
rect 7356 28858 7412 28860
rect 7436 28858 7492 28860
rect 7516 28858 7572 28860
rect 7596 28858 7652 28860
rect 7356 28806 7402 28858
rect 7402 28806 7412 28858
rect 7436 28806 7466 28858
rect 7466 28806 7478 28858
rect 7478 28806 7492 28858
rect 7516 28806 7530 28858
rect 7530 28806 7542 28858
rect 7542 28806 7572 28858
rect 7596 28806 7606 28858
rect 7606 28806 7652 28858
rect 7356 28804 7412 28806
rect 7436 28804 7492 28806
rect 7516 28804 7572 28806
rect 7596 28804 7652 28806
rect 7356 27770 7412 27772
rect 7436 27770 7492 27772
rect 7516 27770 7572 27772
rect 7596 27770 7652 27772
rect 7356 27718 7402 27770
rect 7402 27718 7412 27770
rect 7436 27718 7466 27770
rect 7466 27718 7478 27770
rect 7478 27718 7492 27770
rect 7516 27718 7530 27770
rect 7530 27718 7542 27770
rect 7542 27718 7572 27770
rect 7596 27718 7606 27770
rect 7606 27718 7652 27770
rect 7356 27716 7412 27718
rect 7436 27716 7492 27718
rect 7516 27716 7572 27718
rect 7596 27716 7652 27718
rect 8016 41370 8072 41372
rect 8096 41370 8152 41372
rect 8176 41370 8232 41372
rect 8256 41370 8312 41372
rect 8016 41318 8062 41370
rect 8062 41318 8072 41370
rect 8096 41318 8126 41370
rect 8126 41318 8138 41370
rect 8138 41318 8152 41370
rect 8176 41318 8190 41370
rect 8190 41318 8202 41370
rect 8202 41318 8232 41370
rect 8256 41318 8266 41370
rect 8266 41318 8312 41370
rect 8016 41316 8072 41318
rect 8096 41316 8152 41318
rect 8176 41316 8232 41318
rect 8256 41316 8312 41318
rect 8390 40568 8446 40624
rect 8016 40282 8072 40284
rect 8096 40282 8152 40284
rect 8176 40282 8232 40284
rect 8256 40282 8312 40284
rect 8016 40230 8062 40282
rect 8062 40230 8072 40282
rect 8096 40230 8126 40282
rect 8126 40230 8138 40282
rect 8138 40230 8152 40282
rect 8176 40230 8190 40282
rect 8190 40230 8202 40282
rect 8202 40230 8232 40282
rect 8256 40230 8266 40282
rect 8266 40230 8312 40282
rect 8016 40228 8072 40230
rect 8096 40228 8152 40230
rect 8176 40228 8232 40230
rect 8256 40228 8312 40230
rect 8390 39208 8446 39264
rect 8016 39194 8072 39196
rect 8096 39194 8152 39196
rect 8176 39194 8232 39196
rect 8256 39194 8312 39196
rect 8016 39142 8062 39194
rect 8062 39142 8072 39194
rect 8096 39142 8126 39194
rect 8126 39142 8138 39194
rect 8138 39142 8152 39194
rect 8176 39142 8190 39194
rect 8190 39142 8202 39194
rect 8202 39142 8232 39194
rect 8256 39142 8266 39194
rect 8266 39142 8312 39194
rect 8016 39140 8072 39142
rect 8096 39140 8152 39142
rect 8176 39140 8232 39142
rect 8256 39140 8312 39142
rect 8016 38106 8072 38108
rect 8096 38106 8152 38108
rect 8176 38106 8232 38108
rect 8256 38106 8312 38108
rect 8016 38054 8062 38106
rect 8062 38054 8072 38106
rect 8096 38054 8126 38106
rect 8126 38054 8138 38106
rect 8138 38054 8152 38106
rect 8176 38054 8190 38106
rect 8190 38054 8202 38106
rect 8202 38054 8232 38106
rect 8256 38054 8266 38106
rect 8266 38054 8312 38106
rect 8016 38052 8072 38054
rect 8096 38052 8152 38054
rect 8176 38052 8232 38054
rect 8256 38052 8312 38054
rect 8390 37848 8446 37904
rect 8016 37018 8072 37020
rect 8096 37018 8152 37020
rect 8176 37018 8232 37020
rect 8256 37018 8312 37020
rect 8016 36966 8062 37018
rect 8062 36966 8072 37018
rect 8096 36966 8126 37018
rect 8126 36966 8138 37018
rect 8138 36966 8152 37018
rect 8176 36966 8190 37018
rect 8190 36966 8202 37018
rect 8202 36966 8232 37018
rect 8256 36966 8266 37018
rect 8266 36966 8312 37018
rect 8016 36964 8072 36966
rect 8096 36964 8152 36966
rect 8176 36964 8232 36966
rect 8256 36964 8312 36966
rect 8390 36488 8446 36544
rect 8016 35930 8072 35932
rect 8096 35930 8152 35932
rect 8176 35930 8232 35932
rect 8256 35930 8312 35932
rect 8016 35878 8062 35930
rect 8062 35878 8072 35930
rect 8096 35878 8126 35930
rect 8126 35878 8138 35930
rect 8138 35878 8152 35930
rect 8176 35878 8190 35930
rect 8190 35878 8202 35930
rect 8202 35878 8232 35930
rect 8256 35878 8266 35930
rect 8266 35878 8312 35930
rect 8016 35876 8072 35878
rect 8096 35876 8152 35878
rect 8176 35876 8232 35878
rect 8256 35876 8312 35878
rect 8390 35128 8446 35184
rect 8016 34842 8072 34844
rect 8096 34842 8152 34844
rect 8176 34842 8232 34844
rect 8256 34842 8312 34844
rect 8016 34790 8062 34842
rect 8062 34790 8072 34842
rect 8096 34790 8126 34842
rect 8126 34790 8138 34842
rect 8138 34790 8152 34842
rect 8176 34790 8190 34842
rect 8190 34790 8202 34842
rect 8202 34790 8232 34842
rect 8256 34790 8266 34842
rect 8266 34790 8312 34842
rect 8016 34788 8072 34790
rect 8096 34788 8152 34790
rect 8176 34788 8232 34790
rect 8256 34788 8312 34790
rect 8016 33754 8072 33756
rect 8096 33754 8152 33756
rect 8176 33754 8232 33756
rect 8256 33754 8312 33756
rect 8016 33702 8062 33754
rect 8062 33702 8072 33754
rect 8096 33702 8126 33754
rect 8126 33702 8138 33754
rect 8138 33702 8152 33754
rect 8176 33702 8190 33754
rect 8190 33702 8202 33754
rect 8202 33702 8232 33754
rect 8256 33702 8266 33754
rect 8266 33702 8312 33754
rect 8016 33700 8072 33702
rect 8096 33700 8152 33702
rect 8176 33700 8232 33702
rect 8256 33700 8312 33702
rect 8016 32666 8072 32668
rect 8096 32666 8152 32668
rect 8176 32666 8232 32668
rect 8256 32666 8312 32668
rect 8016 32614 8062 32666
rect 8062 32614 8072 32666
rect 8096 32614 8126 32666
rect 8126 32614 8138 32666
rect 8138 32614 8152 32666
rect 8176 32614 8190 32666
rect 8190 32614 8202 32666
rect 8202 32614 8232 32666
rect 8256 32614 8266 32666
rect 8266 32614 8312 32666
rect 8016 32612 8072 32614
rect 8096 32612 8152 32614
rect 8176 32612 8232 32614
rect 8256 32612 8312 32614
rect 8666 32408 8722 32464
rect 8016 31578 8072 31580
rect 8096 31578 8152 31580
rect 8176 31578 8232 31580
rect 8256 31578 8312 31580
rect 8016 31526 8062 31578
rect 8062 31526 8072 31578
rect 8096 31526 8126 31578
rect 8126 31526 8138 31578
rect 8138 31526 8152 31578
rect 8176 31526 8190 31578
rect 8190 31526 8202 31578
rect 8202 31526 8232 31578
rect 8256 31526 8266 31578
rect 8266 31526 8312 31578
rect 8016 31524 8072 31526
rect 8096 31524 8152 31526
rect 8176 31524 8232 31526
rect 8256 31524 8312 31526
rect 8390 31048 8446 31104
rect 8016 30490 8072 30492
rect 8096 30490 8152 30492
rect 8176 30490 8232 30492
rect 8256 30490 8312 30492
rect 8016 30438 8062 30490
rect 8062 30438 8072 30490
rect 8096 30438 8126 30490
rect 8126 30438 8138 30490
rect 8138 30438 8152 30490
rect 8176 30438 8190 30490
rect 8190 30438 8202 30490
rect 8202 30438 8232 30490
rect 8256 30438 8266 30490
rect 8266 30438 8312 30490
rect 8016 30436 8072 30438
rect 8096 30436 8152 30438
rect 8176 30436 8232 30438
rect 8256 30436 8312 30438
rect 8390 29688 8446 29744
rect 8016 29402 8072 29404
rect 8096 29402 8152 29404
rect 8176 29402 8232 29404
rect 8256 29402 8312 29404
rect 8016 29350 8062 29402
rect 8062 29350 8072 29402
rect 8096 29350 8126 29402
rect 8126 29350 8138 29402
rect 8138 29350 8152 29402
rect 8176 29350 8190 29402
rect 8190 29350 8202 29402
rect 8202 29350 8232 29402
rect 8256 29350 8266 29402
rect 8266 29350 8312 29402
rect 8016 29348 8072 29350
rect 8096 29348 8152 29350
rect 8176 29348 8232 29350
rect 8256 29348 8312 29350
rect 8390 28328 8446 28384
rect 8016 28314 8072 28316
rect 8096 28314 8152 28316
rect 8176 28314 8232 28316
rect 8256 28314 8312 28316
rect 8016 28262 8062 28314
rect 8062 28262 8072 28314
rect 8096 28262 8126 28314
rect 8126 28262 8138 28314
rect 8138 28262 8152 28314
rect 8176 28262 8190 28314
rect 8190 28262 8202 28314
rect 8202 28262 8232 28314
rect 8256 28262 8266 28314
rect 8266 28262 8312 28314
rect 8016 28260 8072 28262
rect 8096 28260 8152 28262
rect 8176 28260 8232 28262
rect 8256 28260 8312 28262
rect 7356 26682 7412 26684
rect 7436 26682 7492 26684
rect 7516 26682 7572 26684
rect 7596 26682 7652 26684
rect 7356 26630 7402 26682
rect 7402 26630 7412 26682
rect 7436 26630 7466 26682
rect 7466 26630 7478 26682
rect 7478 26630 7492 26682
rect 7516 26630 7530 26682
rect 7530 26630 7542 26682
rect 7542 26630 7572 26682
rect 7596 26630 7606 26682
rect 7606 26630 7652 26682
rect 7356 26628 7412 26630
rect 7436 26628 7492 26630
rect 7516 26628 7572 26630
rect 7596 26628 7652 26630
rect 7746 25608 7802 25664
rect 7356 25594 7412 25596
rect 7436 25594 7492 25596
rect 7516 25594 7572 25596
rect 7596 25594 7652 25596
rect 7356 25542 7402 25594
rect 7402 25542 7412 25594
rect 7436 25542 7466 25594
rect 7466 25542 7478 25594
rect 7478 25542 7492 25594
rect 7516 25542 7530 25594
rect 7530 25542 7542 25594
rect 7542 25542 7572 25594
rect 7596 25542 7606 25594
rect 7606 25542 7652 25594
rect 7356 25540 7412 25542
rect 7436 25540 7492 25542
rect 7516 25540 7572 25542
rect 7596 25540 7652 25542
rect 8016 27226 8072 27228
rect 8096 27226 8152 27228
rect 8176 27226 8232 27228
rect 8256 27226 8312 27228
rect 8016 27174 8062 27226
rect 8062 27174 8072 27226
rect 8096 27174 8126 27226
rect 8126 27174 8138 27226
rect 8138 27174 8152 27226
rect 8176 27174 8190 27226
rect 8190 27174 8202 27226
rect 8202 27174 8232 27226
rect 8256 27174 8266 27226
rect 8266 27174 8312 27226
rect 8016 27172 8072 27174
rect 8096 27172 8152 27174
rect 8176 27172 8232 27174
rect 8256 27172 8312 27174
rect 8850 26968 8906 27024
rect 8016 26138 8072 26140
rect 8096 26138 8152 26140
rect 8176 26138 8232 26140
rect 8256 26138 8312 26140
rect 8016 26086 8062 26138
rect 8062 26086 8072 26138
rect 8096 26086 8126 26138
rect 8126 26086 8138 26138
rect 8138 26086 8152 26138
rect 8176 26086 8190 26138
rect 8190 26086 8202 26138
rect 8202 26086 8232 26138
rect 8256 26086 8266 26138
rect 8266 26086 8312 26138
rect 8016 26084 8072 26086
rect 8096 26084 8152 26086
rect 8176 26084 8232 26086
rect 8256 26084 8312 26086
rect 8016 25050 8072 25052
rect 8096 25050 8152 25052
rect 8176 25050 8232 25052
rect 8256 25050 8312 25052
rect 8016 24998 8062 25050
rect 8062 24998 8072 25050
rect 8096 24998 8126 25050
rect 8126 24998 8138 25050
rect 8138 24998 8152 25050
rect 8176 24998 8190 25050
rect 8190 24998 8202 25050
rect 8202 24998 8232 25050
rect 8256 24998 8266 25050
rect 8266 24998 8312 25050
rect 8016 24996 8072 24998
rect 8096 24996 8152 24998
rect 8176 24996 8232 24998
rect 8256 24996 8312 24998
rect 7356 24506 7412 24508
rect 7436 24506 7492 24508
rect 7516 24506 7572 24508
rect 7596 24506 7652 24508
rect 7356 24454 7402 24506
rect 7402 24454 7412 24506
rect 7436 24454 7466 24506
rect 7466 24454 7478 24506
rect 7478 24454 7492 24506
rect 7516 24454 7530 24506
rect 7530 24454 7542 24506
rect 7542 24454 7572 24506
rect 7596 24454 7606 24506
rect 7606 24454 7652 24506
rect 7356 24452 7412 24454
rect 7436 24452 7492 24454
rect 7516 24452 7572 24454
rect 7596 24452 7652 24454
rect 7378 24248 7434 24304
rect 7356 23418 7412 23420
rect 7436 23418 7492 23420
rect 7516 23418 7572 23420
rect 7596 23418 7652 23420
rect 7356 23366 7402 23418
rect 7402 23366 7412 23418
rect 7436 23366 7466 23418
rect 7466 23366 7478 23418
rect 7478 23366 7492 23418
rect 7516 23366 7530 23418
rect 7530 23366 7542 23418
rect 7542 23366 7572 23418
rect 7596 23366 7606 23418
rect 7606 23366 7652 23418
rect 7356 23364 7412 23366
rect 7436 23364 7492 23366
rect 7516 23364 7572 23366
rect 7596 23364 7652 23366
rect 8016 23962 8072 23964
rect 8096 23962 8152 23964
rect 8176 23962 8232 23964
rect 8256 23962 8312 23964
rect 8016 23910 8062 23962
rect 8062 23910 8072 23962
rect 8096 23910 8126 23962
rect 8126 23910 8138 23962
rect 8138 23910 8152 23962
rect 8176 23910 8190 23962
rect 8190 23910 8202 23962
rect 8202 23910 8232 23962
rect 8256 23910 8266 23962
rect 8266 23910 8312 23962
rect 8016 23908 8072 23910
rect 8096 23908 8152 23910
rect 8176 23908 8232 23910
rect 8256 23908 8312 23910
rect 8390 22888 8446 22944
rect 8016 22874 8072 22876
rect 8096 22874 8152 22876
rect 8176 22874 8232 22876
rect 8256 22874 8312 22876
rect 8016 22822 8062 22874
rect 8062 22822 8072 22874
rect 8096 22822 8126 22874
rect 8126 22822 8138 22874
rect 8138 22822 8152 22874
rect 8176 22822 8190 22874
rect 8190 22822 8202 22874
rect 8202 22822 8232 22874
rect 8256 22822 8266 22874
rect 8266 22822 8312 22874
rect 8016 22820 8072 22822
rect 8096 22820 8152 22822
rect 8176 22820 8232 22822
rect 8256 22820 8312 22822
rect 7356 22330 7412 22332
rect 7436 22330 7492 22332
rect 7516 22330 7572 22332
rect 7596 22330 7652 22332
rect 7356 22278 7402 22330
rect 7402 22278 7412 22330
rect 7436 22278 7466 22330
rect 7466 22278 7478 22330
rect 7478 22278 7492 22330
rect 7516 22278 7530 22330
rect 7530 22278 7542 22330
rect 7542 22278 7572 22330
rect 7596 22278 7606 22330
rect 7606 22278 7652 22330
rect 7356 22276 7412 22278
rect 7436 22276 7492 22278
rect 7516 22276 7572 22278
rect 7596 22276 7652 22278
rect 8016 21786 8072 21788
rect 8096 21786 8152 21788
rect 8176 21786 8232 21788
rect 8256 21786 8312 21788
rect 8016 21734 8062 21786
rect 8062 21734 8072 21786
rect 8096 21734 8126 21786
rect 8126 21734 8138 21786
rect 8138 21734 8152 21786
rect 8176 21734 8190 21786
rect 8190 21734 8202 21786
rect 8202 21734 8232 21786
rect 8256 21734 8266 21786
rect 8266 21734 8312 21786
rect 8016 21732 8072 21734
rect 8096 21732 8152 21734
rect 8176 21732 8232 21734
rect 8256 21732 8312 21734
rect 8298 21564 8300 21584
rect 8300 21564 8352 21584
rect 8352 21564 8354 21584
rect 8298 21528 8354 21564
rect 7356 21242 7412 21244
rect 7436 21242 7492 21244
rect 7516 21242 7572 21244
rect 7596 21242 7652 21244
rect 7356 21190 7402 21242
rect 7402 21190 7412 21242
rect 7436 21190 7466 21242
rect 7466 21190 7478 21242
rect 7478 21190 7492 21242
rect 7516 21190 7530 21242
rect 7530 21190 7542 21242
rect 7542 21190 7572 21242
rect 7596 21190 7606 21242
rect 7606 21190 7652 21242
rect 7356 21188 7412 21190
rect 7436 21188 7492 21190
rect 7516 21188 7572 21190
rect 7596 21188 7652 21190
rect 8016 20698 8072 20700
rect 8096 20698 8152 20700
rect 8176 20698 8232 20700
rect 8256 20698 8312 20700
rect 8016 20646 8062 20698
rect 8062 20646 8072 20698
rect 8096 20646 8126 20698
rect 8126 20646 8138 20698
rect 8138 20646 8152 20698
rect 8176 20646 8190 20698
rect 8190 20646 8202 20698
rect 8202 20646 8232 20698
rect 8256 20646 8266 20698
rect 8266 20646 8312 20698
rect 8016 20644 8072 20646
rect 8096 20644 8152 20646
rect 8176 20644 8232 20646
rect 8256 20644 8312 20646
rect 7356 20154 7412 20156
rect 7436 20154 7492 20156
rect 7516 20154 7572 20156
rect 7596 20154 7652 20156
rect 7356 20102 7402 20154
rect 7402 20102 7412 20154
rect 7436 20102 7466 20154
rect 7466 20102 7478 20154
rect 7478 20102 7492 20154
rect 7516 20102 7530 20154
rect 7530 20102 7542 20154
rect 7542 20102 7572 20154
rect 7596 20102 7606 20154
rect 7606 20102 7652 20154
rect 7356 20100 7412 20102
rect 7436 20100 7492 20102
rect 7516 20100 7572 20102
rect 7596 20100 7652 20102
rect 7356 19066 7412 19068
rect 7436 19066 7492 19068
rect 7516 19066 7572 19068
rect 7596 19066 7652 19068
rect 7356 19014 7402 19066
rect 7402 19014 7412 19066
rect 7436 19014 7466 19066
rect 7466 19014 7478 19066
rect 7478 19014 7492 19066
rect 7516 19014 7530 19066
rect 7530 19014 7542 19066
rect 7542 19014 7572 19066
rect 7596 19014 7606 19066
rect 7606 19014 7652 19066
rect 7356 19012 7412 19014
rect 7436 19012 7492 19014
rect 7516 19012 7572 19014
rect 7596 19012 7652 19014
rect 8298 20168 8354 20224
rect 8016 19610 8072 19612
rect 8096 19610 8152 19612
rect 8176 19610 8232 19612
rect 8256 19610 8312 19612
rect 8016 19558 8062 19610
rect 8062 19558 8072 19610
rect 8096 19558 8126 19610
rect 8126 19558 8138 19610
rect 8138 19558 8152 19610
rect 8176 19558 8190 19610
rect 8190 19558 8202 19610
rect 8202 19558 8232 19610
rect 8256 19558 8266 19610
rect 8266 19558 8312 19610
rect 8016 19556 8072 19558
rect 8096 19556 8152 19558
rect 8176 19556 8232 19558
rect 8256 19556 8312 19558
rect 8206 18808 8262 18864
rect 8016 18522 8072 18524
rect 8096 18522 8152 18524
rect 8176 18522 8232 18524
rect 8256 18522 8312 18524
rect 8016 18470 8062 18522
rect 8062 18470 8072 18522
rect 8096 18470 8126 18522
rect 8126 18470 8138 18522
rect 8138 18470 8152 18522
rect 8176 18470 8190 18522
rect 8190 18470 8202 18522
rect 8202 18470 8232 18522
rect 8256 18470 8266 18522
rect 8266 18470 8312 18522
rect 8016 18468 8072 18470
rect 8096 18468 8152 18470
rect 8176 18468 8232 18470
rect 8256 18468 8312 18470
rect 7356 17978 7412 17980
rect 7436 17978 7492 17980
rect 7516 17978 7572 17980
rect 7596 17978 7652 17980
rect 7356 17926 7402 17978
rect 7402 17926 7412 17978
rect 7436 17926 7466 17978
rect 7466 17926 7478 17978
rect 7478 17926 7492 17978
rect 7516 17926 7530 17978
rect 7530 17926 7542 17978
rect 7542 17926 7572 17978
rect 7596 17926 7606 17978
rect 7606 17926 7652 17978
rect 7356 17924 7412 17926
rect 7436 17924 7492 17926
rect 7516 17924 7572 17926
rect 7596 17924 7652 17926
rect 2356 12538 2412 12540
rect 2436 12538 2492 12540
rect 2516 12538 2572 12540
rect 2596 12538 2652 12540
rect 2356 12486 2402 12538
rect 2402 12486 2412 12538
rect 2436 12486 2466 12538
rect 2466 12486 2478 12538
rect 2478 12486 2492 12538
rect 2516 12486 2530 12538
rect 2530 12486 2542 12538
rect 2542 12486 2572 12538
rect 2596 12486 2606 12538
rect 2606 12486 2652 12538
rect 2356 12484 2412 12486
rect 2436 12484 2492 12486
rect 2516 12484 2572 12486
rect 2596 12484 2652 12486
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 3176 11994 3232 11996
rect 3256 11994 3312 11996
rect 3016 11942 3062 11994
rect 3062 11942 3072 11994
rect 3096 11942 3126 11994
rect 3126 11942 3138 11994
rect 3138 11942 3152 11994
rect 3176 11942 3190 11994
rect 3190 11942 3202 11994
rect 3202 11942 3232 11994
rect 3256 11942 3266 11994
rect 3266 11942 3312 11994
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 3176 11940 3232 11942
rect 3256 11940 3312 11942
rect 2356 11450 2412 11452
rect 2436 11450 2492 11452
rect 2516 11450 2572 11452
rect 2596 11450 2652 11452
rect 2356 11398 2402 11450
rect 2402 11398 2412 11450
rect 2436 11398 2466 11450
rect 2466 11398 2478 11450
rect 2478 11398 2492 11450
rect 2516 11398 2530 11450
rect 2530 11398 2542 11450
rect 2542 11398 2572 11450
rect 2596 11398 2606 11450
rect 2606 11398 2652 11450
rect 2356 11396 2412 11398
rect 2436 11396 2492 11398
rect 2516 11396 2572 11398
rect 2596 11396 2652 11398
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 3176 10906 3232 10908
rect 3256 10906 3312 10908
rect 3016 10854 3062 10906
rect 3062 10854 3072 10906
rect 3096 10854 3126 10906
rect 3126 10854 3138 10906
rect 3138 10854 3152 10906
rect 3176 10854 3190 10906
rect 3190 10854 3202 10906
rect 3202 10854 3232 10906
rect 3256 10854 3266 10906
rect 3266 10854 3312 10906
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 3176 10852 3232 10854
rect 3256 10852 3312 10854
rect 2356 10362 2412 10364
rect 2436 10362 2492 10364
rect 2516 10362 2572 10364
rect 2596 10362 2652 10364
rect 2356 10310 2402 10362
rect 2402 10310 2412 10362
rect 2436 10310 2466 10362
rect 2466 10310 2478 10362
rect 2478 10310 2492 10362
rect 2516 10310 2530 10362
rect 2530 10310 2542 10362
rect 2542 10310 2572 10362
rect 2596 10310 2606 10362
rect 2606 10310 2652 10362
rect 2356 10308 2412 10310
rect 2436 10308 2492 10310
rect 2516 10308 2572 10310
rect 2596 10308 2652 10310
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 3176 9818 3232 9820
rect 3256 9818 3312 9820
rect 3016 9766 3062 9818
rect 3062 9766 3072 9818
rect 3096 9766 3126 9818
rect 3126 9766 3138 9818
rect 3138 9766 3152 9818
rect 3176 9766 3190 9818
rect 3190 9766 3202 9818
rect 3202 9766 3232 9818
rect 3256 9766 3266 9818
rect 3266 9766 3312 9818
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 3176 9764 3232 9766
rect 3256 9764 3312 9766
rect 2356 9274 2412 9276
rect 2436 9274 2492 9276
rect 2516 9274 2572 9276
rect 2596 9274 2652 9276
rect 2356 9222 2402 9274
rect 2402 9222 2412 9274
rect 2436 9222 2466 9274
rect 2466 9222 2478 9274
rect 2478 9222 2492 9274
rect 2516 9222 2530 9274
rect 2530 9222 2542 9274
rect 2542 9222 2572 9274
rect 2596 9222 2606 9274
rect 2606 9222 2652 9274
rect 2356 9220 2412 9222
rect 2436 9220 2492 9222
rect 2516 9220 2572 9222
rect 2596 9220 2652 9222
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 2356 8186 2412 8188
rect 2436 8186 2492 8188
rect 2516 8186 2572 8188
rect 2596 8186 2652 8188
rect 2356 8134 2402 8186
rect 2402 8134 2412 8186
rect 2436 8134 2466 8186
rect 2466 8134 2478 8186
rect 2478 8134 2492 8186
rect 2516 8134 2530 8186
rect 2530 8134 2542 8186
rect 2542 8134 2572 8186
rect 2596 8134 2606 8186
rect 2606 8134 2652 8186
rect 2356 8132 2412 8134
rect 2436 8132 2492 8134
rect 2516 8132 2572 8134
rect 2596 8132 2652 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 2356 7098 2412 7100
rect 2436 7098 2492 7100
rect 2516 7098 2572 7100
rect 2596 7098 2652 7100
rect 2356 7046 2402 7098
rect 2402 7046 2412 7098
rect 2436 7046 2466 7098
rect 2466 7046 2478 7098
rect 2478 7046 2492 7098
rect 2516 7046 2530 7098
rect 2530 7046 2542 7098
rect 2542 7046 2572 7098
rect 2596 7046 2606 7098
rect 2606 7046 2652 7098
rect 2356 7044 2412 7046
rect 2436 7044 2492 7046
rect 2516 7044 2572 7046
rect 2596 7044 2652 7046
rect 8016 17434 8072 17436
rect 8096 17434 8152 17436
rect 8176 17434 8232 17436
rect 8256 17434 8312 17436
rect 8016 17382 8062 17434
rect 8062 17382 8072 17434
rect 8096 17382 8126 17434
rect 8126 17382 8138 17434
rect 8138 17382 8152 17434
rect 8176 17382 8190 17434
rect 8190 17382 8202 17434
rect 8202 17382 8232 17434
rect 8256 17382 8266 17434
rect 8266 17382 8312 17434
rect 8016 17380 8072 17382
rect 8096 17380 8152 17382
rect 8176 17380 8232 17382
rect 8256 17380 8312 17382
rect 8482 17448 8538 17504
rect 7356 16890 7412 16892
rect 7436 16890 7492 16892
rect 7516 16890 7572 16892
rect 7596 16890 7652 16892
rect 7356 16838 7402 16890
rect 7402 16838 7412 16890
rect 7436 16838 7466 16890
rect 7466 16838 7478 16890
rect 7478 16838 7492 16890
rect 7516 16838 7530 16890
rect 7530 16838 7542 16890
rect 7542 16838 7572 16890
rect 7596 16838 7606 16890
rect 7606 16838 7652 16890
rect 7356 16836 7412 16838
rect 7436 16836 7492 16838
rect 7516 16836 7572 16838
rect 7596 16836 7652 16838
rect 8016 16346 8072 16348
rect 8096 16346 8152 16348
rect 8176 16346 8232 16348
rect 8256 16346 8312 16348
rect 8016 16294 8062 16346
rect 8062 16294 8072 16346
rect 8096 16294 8126 16346
rect 8126 16294 8138 16346
rect 8138 16294 8152 16346
rect 8176 16294 8190 16346
rect 8190 16294 8202 16346
rect 8202 16294 8232 16346
rect 8256 16294 8266 16346
rect 8266 16294 8312 16346
rect 8016 16292 8072 16294
rect 8096 16292 8152 16294
rect 8176 16292 8232 16294
rect 8256 16292 8312 16294
rect 7356 15802 7412 15804
rect 7436 15802 7492 15804
rect 7516 15802 7572 15804
rect 7596 15802 7652 15804
rect 7356 15750 7402 15802
rect 7402 15750 7412 15802
rect 7436 15750 7466 15802
rect 7466 15750 7478 15802
rect 7478 15750 7492 15802
rect 7516 15750 7530 15802
rect 7530 15750 7542 15802
rect 7542 15750 7572 15802
rect 7596 15750 7606 15802
rect 7606 15750 7652 15802
rect 7356 15748 7412 15750
rect 7436 15748 7492 15750
rect 7516 15748 7572 15750
rect 7596 15748 7652 15750
rect 7356 14714 7412 14716
rect 7436 14714 7492 14716
rect 7516 14714 7572 14716
rect 7596 14714 7652 14716
rect 7356 14662 7402 14714
rect 7402 14662 7412 14714
rect 7436 14662 7466 14714
rect 7466 14662 7478 14714
rect 7478 14662 7492 14714
rect 7516 14662 7530 14714
rect 7530 14662 7542 14714
rect 7542 14662 7572 14714
rect 7596 14662 7606 14714
rect 7606 14662 7652 14714
rect 7356 14660 7412 14662
rect 7436 14660 7492 14662
rect 7516 14660 7572 14662
rect 7596 14660 7652 14662
rect 8016 15258 8072 15260
rect 8096 15258 8152 15260
rect 8176 15258 8232 15260
rect 8256 15258 8312 15260
rect 8016 15206 8062 15258
rect 8062 15206 8072 15258
rect 8096 15206 8126 15258
rect 8126 15206 8138 15258
rect 8138 15206 8152 15258
rect 8176 15206 8190 15258
rect 8190 15206 8202 15258
rect 8202 15206 8232 15258
rect 8256 15206 8266 15258
rect 8266 15206 8312 15258
rect 8016 15204 8072 15206
rect 8096 15204 8152 15206
rect 8176 15204 8232 15206
rect 8256 15204 8312 15206
rect 8850 14728 8906 14784
rect 7356 13626 7412 13628
rect 7436 13626 7492 13628
rect 7516 13626 7572 13628
rect 7596 13626 7652 13628
rect 7356 13574 7402 13626
rect 7402 13574 7412 13626
rect 7436 13574 7466 13626
rect 7466 13574 7478 13626
rect 7478 13574 7492 13626
rect 7516 13574 7530 13626
rect 7530 13574 7542 13626
rect 7542 13574 7572 13626
rect 7596 13574 7606 13626
rect 7606 13574 7652 13626
rect 7356 13572 7412 13574
rect 7436 13572 7492 13574
rect 7516 13572 7572 13574
rect 7596 13572 7652 13574
rect 8016 14170 8072 14172
rect 8096 14170 8152 14172
rect 8176 14170 8232 14172
rect 8256 14170 8312 14172
rect 8016 14118 8062 14170
rect 8062 14118 8072 14170
rect 8096 14118 8126 14170
rect 8126 14118 8138 14170
rect 8138 14118 8152 14170
rect 8176 14118 8190 14170
rect 8190 14118 8202 14170
rect 8202 14118 8232 14170
rect 8256 14118 8266 14170
rect 8266 14118 8312 14170
rect 8016 14116 8072 14118
rect 8096 14116 8152 14118
rect 8176 14116 8232 14118
rect 8256 14116 8312 14118
rect 8298 13368 8354 13424
rect 7356 12538 7412 12540
rect 7436 12538 7492 12540
rect 7516 12538 7572 12540
rect 7596 12538 7652 12540
rect 7356 12486 7402 12538
rect 7402 12486 7412 12538
rect 7436 12486 7466 12538
rect 7466 12486 7478 12538
rect 7478 12486 7492 12538
rect 7516 12486 7530 12538
rect 7530 12486 7542 12538
rect 7542 12486 7572 12538
rect 7596 12486 7606 12538
rect 7606 12486 7652 12538
rect 7356 12484 7412 12486
rect 7436 12484 7492 12486
rect 7516 12484 7572 12486
rect 7596 12484 7652 12486
rect 8016 13082 8072 13084
rect 8096 13082 8152 13084
rect 8176 13082 8232 13084
rect 8256 13082 8312 13084
rect 8016 13030 8062 13082
rect 8062 13030 8072 13082
rect 8096 13030 8126 13082
rect 8126 13030 8138 13082
rect 8138 13030 8152 13082
rect 8176 13030 8190 13082
rect 8190 13030 8202 13082
rect 8202 13030 8232 13082
rect 8256 13030 8266 13082
rect 8266 13030 8312 13082
rect 8016 13028 8072 13030
rect 8096 13028 8152 13030
rect 8176 13028 8232 13030
rect 8256 13028 8312 13030
rect 7010 7928 7066 7984
rect 8016 11994 8072 11996
rect 8096 11994 8152 11996
rect 8176 11994 8232 11996
rect 8256 11994 8312 11996
rect 8016 11942 8062 11994
rect 8062 11942 8072 11994
rect 8096 11942 8126 11994
rect 8126 11942 8138 11994
rect 8138 11942 8152 11994
rect 8176 11942 8190 11994
rect 8190 11942 8202 11994
rect 8202 11942 8232 11994
rect 8256 11942 8266 11994
rect 8266 11942 8312 11994
rect 8016 11940 8072 11942
rect 8096 11940 8152 11942
rect 8176 11940 8232 11942
rect 8256 11940 8312 11942
rect 8482 12008 8538 12064
rect 7356 11450 7412 11452
rect 7436 11450 7492 11452
rect 7516 11450 7572 11452
rect 7596 11450 7652 11452
rect 7356 11398 7402 11450
rect 7402 11398 7412 11450
rect 7436 11398 7466 11450
rect 7466 11398 7478 11450
rect 7478 11398 7492 11450
rect 7516 11398 7530 11450
rect 7530 11398 7542 11450
rect 7542 11398 7572 11450
rect 7596 11398 7606 11450
rect 7606 11398 7652 11450
rect 7356 11396 7412 11398
rect 7436 11396 7492 11398
rect 7516 11396 7572 11398
rect 7596 11396 7652 11398
rect 8016 10906 8072 10908
rect 8096 10906 8152 10908
rect 8176 10906 8232 10908
rect 8256 10906 8312 10908
rect 8016 10854 8062 10906
rect 8062 10854 8072 10906
rect 8096 10854 8126 10906
rect 8126 10854 8138 10906
rect 8138 10854 8152 10906
rect 8176 10854 8190 10906
rect 8190 10854 8202 10906
rect 8202 10854 8232 10906
rect 8256 10854 8266 10906
rect 8266 10854 8312 10906
rect 8016 10852 8072 10854
rect 8096 10852 8152 10854
rect 8176 10852 8232 10854
rect 8256 10852 8312 10854
rect 7930 10648 7986 10704
rect 7356 10362 7412 10364
rect 7436 10362 7492 10364
rect 7516 10362 7572 10364
rect 7596 10362 7652 10364
rect 7356 10310 7402 10362
rect 7402 10310 7412 10362
rect 7436 10310 7466 10362
rect 7466 10310 7478 10362
rect 7478 10310 7492 10362
rect 7516 10310 7530 10362
rect 7530 10310 7542 10362
rect 7542 10310 7572 10362
rect 7596 10310 7606 10362
rect 7606 10310 7652 10362
rect 7356 10308 7412 10310
rect 7436 10308 7492 10310
rect 7516 10308 7572 10310
rect 7596 10308 7652 10310
rect 8016 9818 8072 9820
rect 8096 9818 8152 9820
rect 8176 9818 8232 9820
rect 8256 9818 8312 9820
rect 8016 9766 8062 9818
rect 8062 9766 8072 9818
rect 8096 9766 8126 9818
rect 8126 9766 8138 9818
rect 8138 9766 8152 9818
rect 8176 9766 8190 9818
rect 8190 9766 8202 9818
rect 8202 9766 8232 9818
rect 8256 9766 8266 9818
rect 8266 9766 8312 9818
rect 8016 9764 8072 9766
rect 8096 9764 8152 9766
rect 8176 9764 8232 9766
rect 8256 9764 8312 9766
rect 7356 9274 7412 9276
rect 7436 9274 7492 9276
rect 7516 9274 7572 9276
rect 7596 9274 7652 9276
rect 7356 9222 7402 9274
rect 7402 9222 7412 9274
rect 7436 9222 7466 9274
rect 7466 9222 7478 9274
rect 7478 9222 7492 9274
rect 7516 9222 7530 9274
rect 7530 9222 7542 9274
rect 7542 9222 7572 9274
rect 7596 9222 7606 9274
rect 7606 9222 7652 9274
rect 7356 9220 7412 9222
rect 7436 9220 7492 9222
rect 7516 9220 7572 9222
rect 7596 9220 7652 9222
rect 7356 8186 7412 8188
rect 7436 8186 7492 8188
rect 7516 8186 7572 8188
rect 7596 8186 7652 8188
rect 7356 8134 7402 8186
rect 7402 8134 7412 8186
rect 7436 8134 7466 8186
rect 7466 8134 7478 8186
rect 7478 8134 7492 8186
rect 7516 8134 7530 8186
rect 7530 8134 7542 8186
rect 7542 8134 7572 8186
rect 7596 8134 7606 8186
rect 7606 8134 7652 8186
rect 7356 8132 7412 8134
rect 7436 8132 7492 8134
rect 7516 8132 7572 8134
rect 7596 8132 7652 8134
rect 8298 9288 8354 9344
rect 8016 8730 8072 8732
rect 8096 8730 8152 8732
rect 8176 8730 8232 8732
rect 8256 8730 8312 8732
rect 8016 8678 8062 8730
rect 8062 8678 8072 8730
rect 8096 8678 8126 8730
rect 8126 8678 8138 8730
rect 8138 8678 8152 8730
rect 8176 8678 8190 8730
rect 8190 8678 8202 8730
rect 8202 8678 8232 8730
rect 8256 8678 8266 8730
rect 8266 8678 8312 8730
rect 8016 8676 8072 8678
rect 8096 8676 8152 8678
rect 8176 8676 8232 8678
rect 8256 8676 8312 8678
rect 7356 7098 7412 7100
rect 7436 7098 7492 7100
rect 7516 7098 7572 7100
rect 7596 7098 7652 7100
rect 7356 7046 7402 7098
rect 7402 7046 7412 7098
rect 7436 7046 7466 7098
rect 7466 7046 7478 7098
rect 7478 7046 7492 7098
rect 7516 7046 7530 7098
rect 7530 7046 7542 7098
rect 7542 7046 7572 7098
rect 7596 7046 7606 7098
rect 7606 7046 7652 7098
rect 7356 7044 7412 7046
rect 7436 7044 7492 7046
rect 7516 7044 7572 7046
rect 7596 7044 7652 7046
rect 7654 6840 7710 6896
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2356 6010 2412 6012
rect 2436 6010 2492 6012
rect 2516 6010 2572 6012
rect 2596 6010 2652 6012
rect 2356 5958 2402 6010
rect 2402 5958 2412 6010
rect 2436 5958 2466 6010
rect 2466 5958 2478 6010
rect 2478 5958 2492 6010
rect 2516 5958 2530 6010
rect 2530 5958 2542 6010
rect 2542 5958 2572 6010
rect 2596 5958 2606 6010
rect 2606 5958 2652 6010
rect 2356 5956 2412 5958
rect 2436 5956 2492 5958
rect 2516 5956 2572 5958
rect 2596 5956 2652 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2356 4922 2412 4924
rect 2436 4922 2492 4924
rect 2516 4922 2572 4924
rect 2596 4922 2652 4924
rect 2356 4870 2402 4922
rect 2402 4870 2412 4922
rect 2436 4870 2466 4922
rect 2466 4870 2478 4922
rect 2478 4870 2492 4922
rect 2516 4870 2530 4922
rect 2530 4870 2542 4922
rect 2542 4870 2572 4922
rect 2596 4870 2606 4922
rect 2606 4870 2652 4922
rect 2356 4868 2412 4870
rect 2436 4868 2492 4870
rect 2516 4868 2572 4870
rect 2596 4868 2652 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2356 3834 2412 3836
rect 2436 3834 2492 3836
rect 2516 3834 2572 3836
rect 2596 3834 2652 3836
rect 2356 3782 2402 3834
rect 2402 3782 2412 3834
rect 2436 3782 2466 3834
rect 2466 3782 2478 3834
rect 2478 3782 2492 3834
rect 2516 3782 2530 3834
rect 2530 3782 2542 3834
rect 2542 3782 2572 3834
rect 2596 3782 2606 3834
rect 2606 3782 2652 3834
rect 2356 3780 2412 3782
rect 2436 3780 2492 3782
rect 2516 3780 2572 3782
rect 2596 3780 2652 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 2356 2746 2412 2748
rect 2436 2746 2492 2748
rect 2516 2746 2572 2748
rect 2596 2746 2652 2748
rect 2356 2694 2402 2746
rect 2402 2694 2412 2746
rect 2436 2694 2466 2746
rect 2466 2694 2478 2746
rect 2478 2694 2492 2746
rect 2516 2694 2530 2746
rect 2530 2694 2542 2746
rect 2542 2694 2572 2746
rect 2596 2694 2606 2746
rect 2606 2694 2652 2746
rect 2356 2692 2412 2694
rect 2436 2692 2492 2694
rect 2516 2692 2572 2694
rect 2596 2692 2652 2694
rect 7356 6010 7412 6012
rect 7436 6010 7492 6012
rect 7516 6010 7572 6012
rect 7596 6010 7652 6012
rect 7356 5958 7402 6010
rect 7402 5958 7412 6010
rect 7436 5958 7466 6010
rect 7466 5958 7478 6010
rect 7478 5958 7492 6010
rect 7516 5958 7530 6010
rect 7530 5958 7542 6010
rect 7542 5958 7572 6010
rect 7596 5958 7606 6010
rect 7606 5958 7652 6010
rect 7356 5956 7412 5958
rect 7436 5956 7492 5958
rect 7516 5956 7572 5958
rect 7596 5956 7652 5958
rect 7356 4922 7412 4924
rect 7436 4922 7492 4924
rect 7516 4922 7572 4924
rect 7596 4922 7652 4924
rect 7356 4870 7402 4922
rect 7402 4870 7412 4922
rect 7436 4870 7466 4922
rect 7466 4870 7478 4922
rect 7478 4870 7492 4922
rect 7516 4870 7530 4922
rect 7530 4870 7542 4922
rect 7542 4870 7572 4922
rect 7596 4870 7606 4922
rect 7606 4870 7652 4922
rect 7356 4868 7412 4870
rect 7436 4868 7492 4870
rect 7516 4868 7572 4870
rect 7596 4868 7652 4870
rect 7356 3834 7412 3836
rect 7436 3834 7492 3836
rect 7516 3834 7572 3836
rect 7596 3834 7652 3836
rect 7356 3782 7402 3834
rect 7402 3782 7412 3834
rect 7436 3782 7466 3834
rect 7466 3782 7478 3834
rect 7478 3782 7492 3834
rect 7516 3782 7530 3834
rect 7530 3782 7542 3834
rect 7542 3782 7572 3834
rect 7596 3782 7606 3834
rect 7606 3782 7652 3834
rect 7356 3780 7412 3782
rect 7436 3780 7492 3782
rect 7516 3780 7572 3782
rect 7596 3780 7652 3782
rect 7356 2746 7412 2748
rect 7436 2746 7492 2748
rect 7516 2746 7572 2748
rect 7596 2746 7652 2748
rect 7356 2694 7402 2746
rect 7402 2694 7412 2746
rect 7436 2694 7466 2746
rect 7466 2694 7478 2746
rect 7478 2694 7492 2746
rect 7516 2694 7530 2746
rect 7530 2694 7542 2746
rect 7542 2694 7572 2746
rect 7596 2694 7606 2746
rect 7606 2694 7652 2746
rect 7356 2692 7412 2694
rect 7436 2692 7492 2694
rect 7516 2692 7572 2694
rect 7596 2692 7652 2694
rect 6642 2624 6698 2680
rect 8016 7642 8072 7644
rect 8096 7642 8152 7644
rect 8176 7642 8232 7644
rect 8256 7642 8312 7644
rect 8016 7590 8062 7642
rect 8062 7590 8072 7642
rect 8096 7590 8126 7642
rect 8126 7590 8138 7642
rect 8138 7590 8152 7642
rect 8176 7590 8190 7642
rect 8190 7590 8202 7642
rect 8202 7590 8232 7642
rect 8256 7590 8266 7642
rect 8266 7590 8312 7642
rect 8016 7588 8072 7590
rect 8096 7588 8152 7590
rect 8176 7588 8232 7590
rect 8256 7588 8312 7590
rect 8016 6554 8072 6556
rect 8096 6554 8152 6556
rect 8176 6554 8232 6556
rect 8256 6554 8312 6556
rect 8016 6502 8062 6554
rect 8062 6502 8072 6554
rect 8096 6502 8126 6554
rect 8126 6502 8138 6554
rect 8138 6502 8152 6554
rect 8176 6502 8190 6554
rect 8190 6502 8202 6554
rect 8202 6502 8232 6554
rect 8256 6502 8266 6554
rect 8266 6502 8312 6554
rect 8016 6500 8072 6502
rect 8096 6500 8152 6502
rect 8176 6500 8232 6502
rect 8256 6500 8312 6502
rect 8850 6568 8906 6624
rect 8016 5466 8072 5468
rect 8096 5466 8152 5468
rect 8176 5466 8232 5468
rect 8256 5466 8312 5468
rect 8016 5414 8062 5466
rect 8062 5414 8072 5466
rect 8096 5414 8126 5466
rect 8126 5414 8138 5466
rect 8138 5414 8152 5466
rect 8176 5414 8190 5466
rect 8190 5414 8202 5466
rect 8202 5414 8232 5466
rect 8256 5414 8266 5466
rect 8266 5414 8312 5466
rect 8016 5412 8072 5414
rect 8096 5412 8152 5414
rect 8176 5412 8232 5414
rect 8256 5412 8312 5414
rect 8016 4378 8072 4380
rect 8096 4378 8152 4380
rect 8176 4378 8232 4380
rect 8256 4378 8312 4380
rect 8016 4326 8062 4378
rect 8062 4326 8072 4378
rect 8096 4326 8126 4378
rect 8126 4326 8138 4378
rect 8138 4326 8152 4378
rect 8176 4326 8190 4378
rect 8190 4326 8202 4378
rect 8202 4326 8232 4378
rect 8256 4326 8266 4378
rect 8266 4326 8312 4378
rect 8016 4324 8072 4326
rect 8096 4324 8152 4326
rect 8176 4324 8232 4326
rect 8256 4324 8312 4326
rect 8016 3290 8072 3292
rect 8096 3290 8152 3292
rect 8176 3290 8232 3292
rect 8256 3290 8312 3292
rect 8016 3238 8062 3290
rect 8062 3238 8072 3290
rect 8096 3238 8126 3290
rect 8126 3238 8138 3290
rect 8138 3238 8152 3290
rect 8176 3238 8190 3290
rect 8190 3238 8202 3290
rect 8202 3238 8232 3290
rect 8256 3238 8266 3290
rect 8266 3238 8312 3290
rect 8016 3236 8072 3238
rect 8096 3236 8152 3238
rect 8176 3236 8232 3238
rect 8256 3236 8312 3238
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 8016 2202 8072 2204
rect 8096 2202 8152 2204
rect 8176 2202 8232 2204
rect 8256 2202 8312 2204
rect 8016 2150 8062 2202
rect 8062 2150 8072 2202
rect 8096 2150 8126 2202
rect 8126 2150 8138 2202
rect 8138 2150 8152 2202
rect 8176 2150 8190 2202
rect 8190 2150 8202 2202
rect 8202 2150 8232 2202
rect 8256 2150 8266 2202
rect 8266 2150 8312 2202
rect 8016 2148 8072 2150
rect 8096 2148 8152 2150
rect 8176 2148 8232 2150
rect 8256 2148 8312 2150
<< metal3 >>
rect 2346 77824 2662 77825
rect 2346 77760 2352 77824
rect 2416 77760 2432 77824
rect 2496 77760 2512 77824
rect 2576 77760 2592 77824
rect 2656 77760 2662 77824
rect 2346 77759 2662 77760
rect 7346 77824 7662 77825
rect 7346 77760 7352 77824
rect 7416 77760 7432 77824
rect 7496 77760 7512 77824
rect 7576 77760 7592 77824
rect 7656 77760 7662 77824
rect 7346 77759 7662 77760
rect 3006 77280 3322 77281
rect 3006 77216 3012 77280
rect 3076 77216 3092 77280
rect 3156 77216 3172 77280
rect 3236 77216 3252 77280
rect 3316 77216 3322 77280
rect 3006 77215 3322 77216
rect 8006 77280 8322 77281
rect 8006 77216 8012 77280
rect 8076 77216 8092 77280
rect 8156 77216 8172 77280
rect 8236 77216 8252 77280
rect 8316 77216 8322 77280
rect 8006 77215 8322 77216
rect 2346 76736 2662 76737
rect 2346 76672 2352 76736
rect 2416 76672 2432 76736
rect 2496 76672 2512 76736
rect 2576 76672 2592 76736
rect 2656 76672 2662 76736
rect 2346 76671 2662 76672
rect 7346 76736 7662 76737
rect 7346 76672 7352 76736
rect 7416 76672 7432 76736
rect 7496 76672 7512 76736
rect 7576 76672 7592 76736
rect 7656 76672 7662 76736
rect 7346 76671 7662 76672
rect 3006 76192 3322 76193
rect 3006 76128 3012 76192
rect 3076 76128 3092 76192
rect 3156 76128 3172 76192
rect 3236 76128 3252 76192
rect 3316 76128 3322 76192
rect 3006 76127 3322 76128
rect 8006 76192 8322 76193
rect 8006 76128 8012 76192
rect 8076 76128 8092 76192
rect 8156 76128 8172 76192
rect 8236 76128 8252 76192
rect 8316 76128 8322 76192
rect 8006 76127 8322 76128
rect 2346 75648 2662 75649
rect 2346 75584 2352 75648
rect 2416 75584 2432 75648
rect 2496 75584 2512 75648
rect 2576 75584 2592 75648
rect 2656 75584 2662 75648
rect 2346 75583 2662 75584
rect 7346 75648 7662 75649
rect 7346 75584 7352 75648
rect 7416 75584 7432 75648
rect 7496 75584 7512 75648
rect 7576 75584 7592 75648
rect 7656 75584 7662 75648
rect 7346 75583 7662 75584
rect 3006 75104 3322 75105
rect 3006 75040 3012 75104
rect 3076 75040 3092 75104
rect 3156 75040 3172 75104
rect 3236 75040 3252 75104
rect 3316 75040 3322 75104
rect 3006 75039 3322 75040
rect 8006 75104 8322 75105
rect 8006 75040 8012 75104
rect 8076 75040 8092 75104
rect 8156 75040 8172 75104
rect 8236 75040 8252 75104
rect 8316 75040 8322 75104
rect 8006 75039 8322 75040
rect 2346 74560 2662 74561
rect 2346 74496 2352 74560
rect 2416 74496 2432 74560
rect 2496 74496 2512 74560
rect 2576 74496 2592 74560
rect 2656 74496 2662 74560
rect 2346 74495 2662 74496
rect 7346 74560 7662 74561
rect 7346 74496 7352 74560
rect 7416 74496 7432 74560
rect 7496 74496 7512 74560
rect 7576 74496 7592 74560
rect 7656 74496 7662 74560
rect 7346 74495 7662 74496
rect 3006 74016 3322 74017
rect 3006 73952 3012 74016
rect 3076 73952 3092 74016
rect 3156 73952 3172 74016
rect 3236 73952 3252 74016
rect 3316 73952 3322 74016
rect 3006 73951 3322 73952
rect 8006 74016 8322 74017
rect 8006 73952 8012 74016
rect 8076 73952 8092 74016
rect 8156 73952 8172 74016
rect 8236 73952 8252 74016
rect 8316 73952 8322 74016
rect 8006 73951 8322 73952
rect 2346 73472 2662 73473
rect 2346 73408 2352 73472
rect 2416 73408 2432 73472
rect 2496 73408 2512 73472
rect 2576 73408 2592 73472
rect 2656 73408 2662 73472
rect 2346 73407 2662 73408
rect 7346 73472 7662 73473
rect 7346 73408 7352 73472
rect 7416 73408 7432 73472
rect 7496 73408 7512 73472
rect 7576 73408 7592 73472
rect 7656 73408 7662 73472
rect 7346 73407 7662 73408
rect 8385 73266 8451 73269
rect 9200 73266 10000 73296
rect 8385 73264 10000 73266
rect 8385 73208 8390 73264
rect 8446 73208 10000 73264
rect 8385 73206 10000 73208
rect 8385 73203 8451 73206
rect 9200 73176 10000 73206
rect 3006 72928 3322 72929
rect 3006 72864 3012 72928
rect 3076 72864 3092 72928
rect 3156 72864 3172 72928
rect 3236 72864 3252 72928
rect 3316 72864 3322 72928
rect 3006 72863 3322 72864
rect 8006 72928 8322 72929
rect 8006 72864 8012 72928
rect 8076 72864 8092 72928
rect 8156 72864 8172 72928
rect 8236 72864 8252 72928
rect 8316 72864 8322 72928
rect 8006 72863 8322 72864
rect 2346 72384 2662 72385
rect 2346 72320 2352 72384
rect 2416 72320 2432 72384
rect 2496 72320 2512 72384
rect 2576 72320 2592 72384
rect 2656 72320 2662 72384
rect 2346 72319 2662 72320
rect 7346 72384 7662 72385
rect 7346 72320 7352 72384
rect 7416 72320 7432 72384
rect 7496 72320 7512 72384
rect 7576 72320 7592 72384
rect 7656 72320 7662 72384
rect 7346 72319 7662 72320
rect 8477 71906 8543 71909
rect 9200 71906 10000 71936
rect 8477 71904 10000 71906
rect 8477 71848 8482 71904
rect 8538 71848 10000 71904
rect 8477 71846 10000 71848
rect 8477 71843 8543 71846
rect 3006 71840 3322 71841
rect 3006 71776 3012 71840
rect 3076 71776 3092 71840
rect 3156 71776 3172 71840
rect 3236 71776 3252 71840
rect 3316 71776 3322 71840
rect 3006 71775 3322 71776
rect 8006 71840 8322 71841
rect 8006 71776 8012 71840
rect 8076 71776 8092 71840
rect 8156 71776 8172 71840
rect 8236 71776 8252 71840
rect 8316 71776 8322 71840
rect 9200 71816 10000 71846
rect 8006 71775 8322 71776
rect 2346 71296 2662 71297
rect 2346 71232 2352 71296
rect 2416 71232 2432 71296
rect 2496 71232 2512 71296
rect 2576 71232 2592 71296
rect 2656 71232 2662 71296
rect 2346 71231 2662 71232
rect 7346 71296 7662 71297
rect 7346 71232 7352 71296
rect 7416 71232 7432 71296
rect 7496 71232 7512 71296
rect 7576 71232 7592 71296
rect 7656 71232 7662 71296
rect 7346 71231 7662 71232
rect 3006 70752 3322 70753
rect 3006 70688 3012 70752
rect 3076 70688 3092 70752
rect 3156 70688 3172 70752
rect 3236 70688 3252 70752
rect 3316 70688 3322 70752
rect 3006 70687 3322 70688
rect 8006 70752 8322 70753
rect 8006 70688 8012 70752
rect 8076 70688 8092 70752
rect 8156 70688 8172 70752
rect 8236 70688 8252 70752
rect 8316 70688 8322 70752
rect 8006 70687 8322 70688
rect 8385 70546 8451 70549
rect 9200 70546 10000 70576
rect 8385 70544 10000 70546
rect 8385 70488 8390 70544
rect 8446 70488 10000 70544
rect 8385 70486 10000 70488
rect 8385 70483 8451 70486
rect 9200 70456 10000 70486
rect 2346 70208 2662 70209
rect 2346 70144 2352 70208
rect 2416 70144 2432 70208
rect 2496 70144 2512 70208
rect 2576 70144 2592 70208
rect 2656 70144 2662 70208
rect 2346 70143 2662 70144
rect 7346 70208 7662 70209
rect 7346 70144 7352 70208
rect 7416 70144 7432 70208
rect 7496 70144 7512 70208
rect 7576 70144 7592 70208
rect 7656 70144 7662 70208
rect 7346 70143 7662 70144
rect 3006 69664 3322 69665
rect 3006 69600 3012 69664
rect 3076 69600 3092 69664
rect 3156 69600 3172 69664
rect 3236 69600 3252 69664
rect 3316 69600 3322 69664
rect 3006 69599 3322 69600
rect 8006 69664 8322 69665
rect 8006 69600 8012 69664
rect 8076 69600 8092 69664
rect 8156 69600 8172 69664
rect 8236 69600 8252 69664
rect 8316 69600 8322 69664
rect 8006 69599 8322 69600
rect 8385 69186 8451 69189
rect 9200 69186 10000 69216
rect 8385 69184 10000 69186
rect 8385 69128 8390 69184
rect 8446 69128 10000 69184
rect 8385 69126 10000 69128
rect 8385 69123 8451 69126
rect 2346 69120 2662 69121
rect 2346 69056 2352 69120
rect 2416 69056 2432 69120
rect 2496 69056 2512 69120
rect 2576 69056 2592 69120
rect 2656 69056 2662 69120
rect 2346 69055 2662 69056
rect 7346 69120 7662 69121
rect 7346 69056 7352 69120
rect 7416 69056 7432 69120
rect 7496 69056 7512 69120
rect 7576 69056 7592 69120
rect 7656 69056 7662 69120
rect 9200 69096 10000 69126
rect 7346 69055 7662 69056
rect 3006 68576 3322 68577
rect 3006 68512 3012 68576
rect 3076 68512 3092 68576
rect 3156 68512 3172 68576
rect 3236 68512 3252 68576
rect 3316 68512 3322 68576
rect 3006 68511 3322 68512
rect 8006 68576 8322 68577
rect 8006 68512 8012 68576
rect 8076 68512 8092 68576
rect 8156 68512 8172 68576
rect 8236 68512 8252 68576
rect 8316 68512 8322 68576
rect 8006 68511 8322 68512
rect 2346 68032 2662 68033
rect 2346 67968 2352 68032
rect 2416 67968 2432 68032
rect 2496 67968 2512 68032
rect 2576 67968 2592 68032
rect 2656 67968 2662 68032
rect 2346 67967 2662 67968
rect 7346 68032 7662 68033
rect 7346 67968 7352 68032
rect 7416 67968 7432 68032
rect 7496 67968 7512 68032
rect 7576 67968 7592 68032
rect 7656 67968 7662 68032
rect 7346 67967 7662 67968
rect 8385 67826 8451 67829
rect 9200 67826 10000 67856
rect 8385 67824 10000 67826
rect 8385 67768 8390 67824
rect 8446 67768 10000 67824
rect 8385 67766 10000 67768
rect 8385 67763 8451 67766
rect 9200 67736 10000 67766
rect 3006 67488 3322 67489
rect 3006 67424 3012 67488
rect 3076 67424 3092 67488
rect 3156 67424 3172 67488
rect 3236 67424 3252 67488
rect 3316 67424 3322 67488
rect 3006 67423 3322 67424
rect 8006 67488 8322 67489
rect 8006 67424 8012 67488
rect 8076 67424 8092 67488
rect 8156 67424 8172 67488
rect 8236 67424 8252 67488
rect 8316 67424 8322 67488
rect 8006 67423 8322 67424
rect 2346 66944 2662 66945
rect 2346 66880 2352 66944
rect 2416 66880 2432 66944
rect 2496 66880 2512 66944
rect 2576 66880 2592 66944
rect 2656 66880 2662 66944
rect 2346 66879 2662 66880
rect 7346 66944 7662 66945
rect 7346 66880 7352 66944
rect 7416 66880 7432 66944
rect 7496 66880 7512 66944
rect 7576 66880 7592 66944
rect 7656 66880 7662 66944
rect 7346 66879 7662 66880
rect 8385 66466 8451 66469
rect 9200 66466 10000 66496
rect 8385 66464 10000 66466
rect 8385 66408 8390 66464
rect 8446 66408 10000 66464
rect 8385 66406 10000 66408
rect 8385 66403 8451 66406
rect 3006 66400 3322 66401
rect 3006 66336 3012 66400
rect 3076 66336 3092 66400
rect 3156 66336 3172 66400
rect 3236 66336 3252 66400
rect 3316 66336 3322 66400
rect 3006 66335 3322 66336
rect 8006 66400 8322 66401
rect 8006 66336 8012 66400
rect 8076 66336 8092 66400
rect 8156 66336 8172 66400
rect 8236 66336 8252 66400
rect 8316 66336 8322 66400
rect 9200 66376 10000 66406
rect 8006 66335 8322 66336
rect 2346 65856 2662 65857
rect 2346 65792 2352 65856
rect 2416 65792 2432 65856
rect 2496 65792 2512 65856
rect 2576 65792 2592 65856
rect 2656 65792 2662 65856
rect 2346 65791 2662 65792
rect 7346 65856 7662 65857
rect 7346 65792 7352 65856
rect 7416 65792 7432 65856
rect 7496 65792 7512 65856
rect 7576 65792 7592 65856
rect 7656 65792 7662 65856
rect 7346 65791 7662 65792
rect 3006 65312 3322 65313
rect 3006 65248 3012 65312
rect 3076 65248 3092 65312
rect 3156 65248 3172 65312
rect 3236 65248 3252 65312
rect 3316 65248 3322 65312
rect 3006 65247 3322 65248
rect 8006 65312 8322 65313
rect 8006 65248 8012 65312
rect 8076 65248 8092 65312
rect 8156 65248 8172 65312
rect 8236 65248 8252 65312
rect 8316 65248 8322 65312
rect 8006 65247 8322 65248
rect 8385 65106 8451 65109
rect 9200 65106 10000 65136
rect 8385 65104 10000 65106
rect 8385 65048 8390 65104
rect 8446 65048 10000 65104
rect 8385 65046 10000 65048
rect 8385 65043 8451 65046
rect 9200 65016 10000 65046
rect 2346 64768 2662 64769
rect 2346 64704 2352 64768
rect 2416 64704 2432 64768
rect 2496 64704 2512 64768
rect 2576 64704 2592 64768
rect 2656 64704 2662 64768
rect 2346 64703 2662 64704
rect 7346 64768 7662 64769
rect 7346 64704 7352 64768
rect 7416 64704 7432 64768
rect 7496 64704 7512 64768
rect 7576 64704 7592 64768
rect 7656 64704 7662 64768
rect 7346 64703 7662 64704
rect 3006 64224 3322 64225
rect 3006 64160 3012 64224
rect 3076 64160 3092 64224
rect 3156 64160 3172 64224
rect 3236 64160 3252 64224
rect 3316 64160 3322 64224
rect 3006 64159 3322 64160
rect 8006 64224 8322 64225
rect 8006 64160 8012 64224
rect 8076 64160 8092 64224
rect 8156 64160 8172 64224
rect 8236 64160 8252 64224
rect 8316 64160 8322 64224
rect 8006 64159 8322 64160
rect 8477 63746 8543 63749
rect 9200 63746 10000 63776
rect 8477 63744 10000 63746
rect 8477 63688 8482 63744
rect 8538 63688 10000 63744
rect 8477 63686 10000 63688
rect 8477 63683 8543 63686
rect 2346 63680 2662 63681
rect 2346 63616 2352 63680
rect 2416 63616 2432 63680
rect 2496 63616 2512 63680
rect 2576 63616 2592 63680
rect 2656 63616 2662 63680
rect 2346 63615 2662 63616
rect 7346 63680 7662 63681
rect 7346 63616 7352 63680
rect 7416 63616 7432 63680
rect 7496 63616 7512 63680
rect 7576 63616 7592 63680
rect 7656 63616 7662 63680
rect 9200 63656 10000 63686
rect 7346 63615 7662 63616
rect 3006 63136 3322 63137
rect 3006 63072 3012 63136
rect 3076 63072 3092 63136
rect 3156 63072 3172 63136
rect 3236 63072 3252 63136
rect 3316 63072 3322 63136
rect 3006 63071 3322 63072
rect 8006 63136 8322 63137
rect 8006 63072 8012 63136
rect 8076 63072 8092 63136
rect 8156 63072 8172 63136
rect 8236 63072 8252 63136
rect 8316 63072 8322 63136
rect 8006 63071 8322 63072
rect 2346 62592 2662 62593
rect 2346 62528 2352 62592
rect 2416 62528 2432 62592
rect 2496 62528 2512 62592
rect 2576 62528 2592 62592
rect 2656 62528 2662 62592
rect 2346 62527 2662 62528
rect 7346 62592 7662 62593
rect 7346 62528 7352 62592
rect 7416 62528 7432 62592
rect 7496 62528 7512 62592
rect 7576 62528 7592 62592
rect 7656 62528 7662 62592
rect 7346 62527 7662 62528
rect 8385 62386 8451 62389
rect 9200 62386 10000 62416
rect 8385 62384 10000 62386
rect 8385 62328 8390 62384
rect 8446 62328 10000 62384
rect 8385 62326 10000 62328
rect 8385 62323 8451 62326
rect 9200 62296 10000 62326
rect 3006 62048 3322 62049
rect 3006 61984 3012 62048
rect 3076 61984 3092 62048
rect 3156 61984 3172 62048
rect 3236 61984 3252 62048
rect 3316 61984 3322 62048
rect 3006 61983 3322 61984
rect 8006 62048 8322 62049
rect 8006 61984 8012 62048
rect 8076 61984 8092 62048
rect 8156 61984 8172 62048
rect 8236 61984 8252 62048
rect 8316 61984 8322 62048
rect 8006 61983 8322 61984
rect 2346 61504 2662 61505
rect 2346 61440 2352 61504
rect 2416 61440 2432 61504
rect 2496 61440 2512 61504
rect 2576 61440 2592 61504
rect 2656 61440 2662 61504
rect 2346 61439 2662 61440
rect 7346 61504 7662 61505
rect 7346 61440 7352 61504
rect 7416 61440 7432 61504
rect 7496 61440 7512 61504
rect 7576 61440 7592 61504
rect 7656 61440 7662 61504
rect 7346 61439 7662 61440
rect 6913 61298 6979 61301
rect 6870 61296 6979 61298
rect 6870 61240 6918 61296
rect 6974 61240 6979 61296
rect 6870 61235 6979 61240
rect 3006 60960 3322 60961
rect 3006 60896 3012 60960
rect 3076 60896 3092 60960
rect 3156 60896 3172 60960
rect 3236 60896 3252 60960
rect 3316 60896 3322 60960
rect 3006 60895 3322 60896
rect 6870 60618 6930 61235
rect 8385 61026 8451 61029
rect 9200 61026 10000 61056
rect 8385 61024 10000 61026
rect 8385 60968 8390 61024
rect 8446 60968 10000 61024
rect 8385 60966 10000 60968
rect 8385 60963 8451 60966
rect 8006 60960 8322 60961
rect 8006 60896 8012 60960
rect 8076 60896 8092 60960
rect 8156 60896 8172 60960
rect 8236 60896 8252 60960
rect 8316 60896 8322 60960
rect 9200 60936 10000 60966
rect 8006 60895 8322 60896
rect 7833 60618 7899 60621
rect 6870 60616 7899 60618
rect 6870 60560 7838 60616
rect 7894 60560 7899 60616
rect 6870 60558 7899 60560
rect 7833 60555 7899 60558
rect 2346 60416 2662 60417
rect 2346 60352 2352 60416
rect 2416 60352 2432 60416
rect 2496 60352 2512 60416
rect 2576 60352 2592 60416
rect 2656 60352 2662 60416
rect 2346 60351 2662 60352
rect 7346 60416 7662 60417
rect 7346 60352 7352 60416
rect 7416 60352 7432 60416
rect 7496 60352 7512 60416
rect 7576 60352 7592 60416
rect 7656 60352 7662 60416
rect 7346 60351 7662 60352
rect 3006 59872 3322 59873
rect 3006 59808 3012 59872
rect 3076 59808 3092 59872
rect 3156 59808 3172 59872
rect 3236 59808 3252 59872
rect 3316 59808 3322 59872
rect 3006 59807 3322 59808
rect 8006 59872 8322 59873
rect 8006 59808 8012 59872
rect 8076 59808 8092 59872
rect 8156 59808 8172 59872
rect 8236 59808 8252 59872
rect 8316 59808 8322 59872
rect 8006 59807 8322 59808
rect 8385 59666 8451 59669
rect 9200 59666 10000 59696
rect 8385 59664 10000 59666
rect 8385 59608 8390 59664
rect 8446 59608 10000 59664
rect 8385 59606 10000 59608
rect 8385 59603 8451 59606
rect 9200 59576 10000 59606
rect 2346 59328 2662 59329
rect 2346 59264 2352 59328
rect 2416 59264 2432 59328
rect 2496 59264 2512 59328
rect 2576 59264 2592 59328
rect 2656 59264 2662 59328
rect 2346 59263 2662 59264
rect 7346 59328 7662 59329
rect 7346 59264 7352 59328
rect 7416 59264 7432 59328
rect 7496 59264 7512 59328
rect 7576 59264 7592 59328
rect 7656 59264 7662 59328
rect 7346 59263 7662 59264
rect 3006 58784 3322 58785
rect 3006 58720 3012 58784
rect 3076 58720 3092 58784
rect 3156 58720 3172 58784
rect 3236 58720 3252 58784
rect 3316 58720 3322 58784
rect 3006 58719 3322 58720
rect 8006 58784 8322 58785
rect 8006 58720 8012 58784
rect 8076 58720 8092 58784
rect 8156 58720 8172 58784
rect 8236 58720 8252 58784
rect 8316 58720 8322 58784
rect 8006 58719 8322 58720
rect 8477 58306 8543 58309
rect 9200 58306 10000 58336
rect 8477 58304 10000 58306
rect 8477 58248 8482 58304
rect 8538 58248 10000 58304
rect 8477 58246 10000 58248
rect 8477 58243 8543 58246
rect 2346 58240 2662 58241
rect 2346 58176 2352 58240
rect 2416 58176 2432 58240
rect 2496 58176 2512 58240
rect 2576 58176 2592 58240
rect 2656 58176 2662 58240
rect 2346 58175 2662 58176
rect 7346 58240 7662 58241
rect 7346 58176 7352 58240
rect 7416 58176 7432 58240
rect 7496 58176 7512 58240
rect 7576 58176 7592 58240
rect 7656 58176 7662 58240
rect 9200 58216 10000 58246
rect 7346 58175 7662 58176
rect 3006 57696 3322 57697
rect 3006 57632 3012 57696
rect 3076 57632 3092 57696
rect 3156 57632 3172 57696
rect 3236 57632 3252 57696
rect 3316 57632 3322 57696
rect 3006 57631 3322 57632
rect 8006 57696 8322 57697
rect 8006 57632 8012 57696
rect 8076 57632 8092 57696
rect 8156 57632 8172 57696
rect 8236 57632 8252 57696
rect 8316 57632 8322 57696
rect 8006 57631 8322 57632
rect 2346 57152 2662 57153
rect 2346 57088 2352 57152
rect 2416 57088 2432 57152
rect 2496 57088 2512 57152
rect 2576 57088 2592 57152
rect 2656 57088 2662 57152
rect 2346 57087 2662 57088
rect 7346 57152 7662 57153
rect 7346 57088 7352 57152
rect 7416 57088 7432 57152
rect 7496 57088 7512 57152
rect 7576 57088 7592 57152
rect 7656 57088 7662 57152
rect 7346 57087 7662 57088
rect 8569 56946 8635 56949
rect 9200 56946 10000 56976
rect 8569 56944 10000 56946
rect 8569 56888 8574 56944
rect 8630 56888 10000 56944
rect 8569 56886 10000 56888
rect 8569 56883 8635 56886
rect 9200 56856 10000 56886
rect 3006 56608 3322 56609
rect 3006 56544 3012 56608
rect 3076 56544 3092 56608
rect 3156 56544 3172 56608
rect 3236 56544 3252 56608
rect 3316 56544 3322 56608
rect 3006 56543 3322 56544
rect 8006 56608 8322 56609
rect 8006 56544 8012 56608
rect 8076 56544 8092 56608
rect 8156 56544 8172 56608
rect 8236 56544 8252 56608
rect 8316 56544 8322 56608
rect 8006 56543 8322 56544
rect 2346 56064 2662 56065
rect 2346 56000 2352 56064
rect 2416 56000 2432 56064
rect 2496 56000 2512 56064
rect 2576 56000 2592 56064
rect 2656 56000 2662 56064
rect 2346 55999 2662 56000
rect 7346 56064 7662 56065
rect 7346 56000 7352 56064
rect 7416 56000 7432 56064
rect 7496 56000 7512 56064
rect 7576 56000 7592 56064
rect 7656 56000 7662 56064
rect 7346 55999 7662 56000
rect 9200 55586 10000 55616
rect 8388 55526 10000 55586
rect 3006 55520 3322 55521
rect 3006 55456 3012 55520
rect 3076 55456 3092 55520
rect 3156 55456 3172 55520
rect 3236 55456 3252 55520
rect 3316 55456 3322 55520
rect 3006 55455 3322 55456
rect 8006 55520 8322 55521
rect 8006 55456 8012 55520
rect 8076 55456 8092 55520
rect 8156 55456 8172 55520
rect 8236 55456 8252 55520
rect 8316 55456 8322 55520
rect 8006 55455 8322 55456
rect 8201 55314 8267 55317
rect 8388 55314 8448 55526
rect 9200 55496 10000 55526
rect 8201 55312 8448 55314
rect 8201 55256 8206 55312
rect 8262 55256 8448 55312
rect 8201 55254 8448 55256
rect 8201 55251 8267 55254
rect 2346 54976 2662 54977
rect 2346 54912 2352 54976
rect 2416 54912 2432 54976
rect 2496 54912 2512 54976
rect 2576 54912 2592 54976
rect 2656 54912 2662 54976
rect 2346 54911 2662 54912
rect 7346 54976 7662 54977
rect 7346 54912 7352 54976
rect 7416 54912 7432 54976
rect 7496 54912 7512 54976
rect 7576 54912 7592 54976
rect 7656 54912 7662 54976
rect 7346 54911 7662 54912
rect 3006 54432 3322 54433
rect 3006 54368 3012 54432
rect 3076 54368 3092 54432
rect 3156 54368 3172 54432
rect 3236 54368 3252 54432
rect 3316 54368 3322 54432
rect 3006 54367 3322 54368
rect 8006 54432 8322 54433
rect 8006 54368 8012 54432
rect 8076 54368 8092 54432
rect 8156 54368 8172 54432
rect 8236 54368 8252 54432
rect 8316 54368 8322 54432
rect 8006 54367 8322 54368
rect 8385 54226 8451 54229
rect 9200 54226 10000 54256
rect 8385 54224 10000 54226
rect 8385 54168 8390 54224
rect 8446 54168 10000 54224
rect 8385 54166 10000 54168
rect 8385 54163 8451 54166
rect 9200 54136 10000 54166
rect 2346 53888 2662 53889
rect 2346 53824 2352 53888
rect 2416 53824 2432 53888
rect 2496 53824 2512 53888
rect 2576 53824 2592 53888
rect 2656 53824 2662 53888
rect 2346 53823 2662 53824
rect 7346 53888 7662 53889
rect 7346 53824 7352 53888
rect 7416 53824 7432 53888
rect 7496 53824 7512 53888
rect 7576 53824 7592 53888
rect 7656 53824 7662 53888
rect 7346 53823 7662 53824
rect 3006 53344 3322 53345
rect 3006 53280 3012 53344
rect 3076 53280 3092 53344
rect 3156 53280 3172 53344
rect 3236 53280 3252 53344
rect 3316 53280 3322 53344
rect 3006 53279 3322 53280
rect 8006 53344 8322 53345
rect 8006 53280 8012 53344
rect 8076 53280 8092 53344
rect 8156 53280 8172 53344
rect 8236 53280 8252 53344
rect 8316 53280 8322 53344
rect 8006 53279 8322 53280
rect 8385 52866 8451 52869
rect 9200 52866 10000 52896
rect 8385 52864 10000 52866
rect 8385 52808 8390 52864
rect 8446 52808 10000 52864
rect 8385 52806 10000 52808
rect 8385 52803 8451 52806
rect 2346 52800 2662 52801
rect 2346 52736 2352 52800
rect 2416 52736 2432 52800
rect 2496 52736 2512 52800
rect 2576 52736 2592 52800
rect 2656 52736 2662 52800
rect 2346 52735 2662 52736
rect 7346 52800 7662 52801
rect 7346 52736 7352 52800
rect 7416 52736 7432 52800
rect 7496 52736 7512 52800
rect 7576 52736 7592 52800
rect 7656 52736 7662 52800
rect 9200 52776 10000 52806
rect 7346 52735 7662 52736
rect 3006 52256 3322 52257
rect 3006 52192 3012 52256
rect 3076 52192 3092 52256
rect 3156 52192 3172 52256
rect 3236 52192 3252 52256
rect 3316 52192 3322 52256
rect 3006 52191 3322 52192
rect 8006 52256 8322 52257
rect 8006 52192 8012 52256
rect 8076 52192 8092 52256
rect 8156 52192 8172 52256
rect 8236 52192 8252 52256
rect 8316 52192 8322 52256
rect 8006 52191 8322 52192
rect 2346 51712 2662 51713
rect 2346 51648 2352 51712
rect 2416 51648 2432 51712
rect 2496 51648 2512 51712
rect 2576 51648 2592 51712
rect 2656 51648 2662 51712
rect 2346 51647 2662 51648
rect 7346 51712 7662 51713
rect 7346 51648 7352 51712
rect 7416 51648 7432 51712
rect 7496 51648 7512 51712
rect 7576 51648 7592 51712
rect 7656 51648 7662 51712
rect 7346 51647 7662 51648
rect 8385 51506 8451 51509
rect 9200 51506 10000 51536
rect 8385 51504 10000 51506
rect 8385 51448 8390 51504
rect 8446 51448 10000 51504
rect 8385 51446 10000 51448
rect 8385 51443 8451 51446
rect 9200 51416 10000 51446
rect 3006 51168 3322 51169
rect 3006 51104 3012 51168
rect 3076 51104 3092 51168
rect 3156 51104 3172 51168
rect 3236 51104 3252 51168
rect 3316 51104 3322 51168
rect 3006 51103 3322 51104
rect 8006 51168 8322 51169
rect 8006 51104 8012 51168
rect 8076 51104 8092 51168
rect 8156 51104 8172 51168
rect 8236 51104 8252 51168
rect 8316 51104 8322 51168
rect 8006 51103 8322 51104
rect 2346 50624 2662 50625
rect 2346 50560 2352 50624
rect 2416 50560 2432 50624
rect 2496 50560 2512 50624
rect 2576 50560 2592 50624
rect 2656 50560 2662 50624
rect 2346 50559 2662 50560
rect 7346 50624 7662 50625
rect 7346 50560 7352 50624
rect 7416 50560 7432 50624
rect 7496 50560 7512 50624
rect 7576 50560 7592 50624
rect 7656 50560 7662 50624
rect 7346 50559 7662 50560
rect 8385 50146 8451 50149
rect 9200 50146 10000 50176
rect 8385 50144 10000 50146
rect 8385 50088 8390 50144
rect 8446 50088 10000 50144
rect 8385 50086 10000 50088
rect 8385 50083 8451 50086
rect 3006 50080 3322 50081
rect 3006 50016 3012 50080
rect 3076 50016 3092 50080
rect 3156 50016 3172 50080
rect 3236 50016 3252 50080
rect 3316 50016 3322 50080
rect 3006 50015 3322 50016
rect 8006 50080 8322 50081
rect 8006 50016 8012 50080
rect 8076 50016 8092 50080
rect 8156 50016 8172 50080
rect 8236 50016 8252 50080
rect 8316 50016 8322 50080
rect 9200 50056 10000 50086
rect 8006 50015 8322 50016
rect 2346 49536 2662 49537
rect 2346 49472 2352 49536
rect 2416 49472 2432 49536
rect 2496 49472 2512 49536
rect 2576 49472 2592 49536
rect 2656 49472 2662 49536
rect 2346 49471 2662 49472
rect 7346 49536 7662 49537
rect 7346 49472 7352 49536
rect 7416 49472 7432 49536
rect 7496 49472 7512 49536
rect 7576 49472 7592 49536
rect 7656 49472 7662 49536
rect 7346 49471 7662 49472
rect 3006 48992 3322 48993
rect 3006 48928 3012 48992
rect 3076 48928 3092 48992
rect 3156 48928 3172 48992
rect 3236 48928 3252 48992
rect 3316 48928 3322 48992
rect 3006 48927 3322 48928
rect 8006 48992 8322 48993
rect 8006 48928 8012 48992
rect 8076 48928 8092 48992
rect 8156 48928 8172 48992
rect 8236 48928 8252 48992
rect 8316 48928 8322 48992
rect 8006 48927 8322 48928
rect 8385 48786 8451 48789
rect 9200 48786 10000 48816
rect 8385 48784 10000 48786
rect 8385 48728 8390 48784
rect 8446 48728 10000 48784
rect 8385 48726 10000 48728
rect 8385 48723 8451 48726
rect 9200 48696 10000 48726
rect 2346 48448 2662 48449
rect 2346 48384 2352 48448
rect 2416 48384 2432 48448
rect 2496 48384 2512 48448
rect 2576 48384 2592 48448
rect 2656 48384 2662 48448
rect 2346 48383 2662 48384
rect 7346 48448 7662 48449
rect 7346 48384 7352 48448
rect 7416 48384 7432 48448
rect 7496 48384 7512 48448
rect 7576 48384 7592 48448
rect 7656 48384 7662 48448
rect 7346 48383 7662 48384
rect 3006 47904 3322 47905
rect 3006 47840 3012 47904
rect 3076 47840 3092 47904
rect 3156 47840 3172 47904
rect 3236 47840 3252 47904
rect 3316 47840 3322 47904
rect 3006 47839 3322 47840
rect 8006 47904 8322 47905
rect 8006 47840 8012 47904
rect 8076 47840 8092 47904
rect 8156 47840 8172 47904
rect 8236 47840 8252 47904
rect 8316 47840 8322 47904
rect 8006 47839 8322 47840
rect 8385 47426 8451 47429
rect 9200 47426 10000 47456
rect 8385 47424 10000 47426
rect 8385 47368 8390 47424
rect 8446 47368 10000 47424
rect 8385 47366 10000 47368
rect 8385 47363 8451 47366
rect 2346 47360 2662 47361
rect 2346 47296 2352 47360
rect 2416 47296 2432 47360
rect 2496 47296 2512 47360
rect 2576 47296 2592 47360
rect 2656 47296 2662 47360
rect 2346 47295 2662 47296
rect 7346 47360 7662 47361
rect 7346 47296 7352 47360
rect 7416 47296 7432 47360
rect 7496 47296 7512 47360
rect 7576 47296 7592 47360
rect 7656 47296 7662 47360
rect 9200 47336 10000 47366
rect 7346 47295 7662 47296
rect 3006 46816 3322 46817
rect 3006 46752 3012 46816
rect 3076 46752 3092 46816
rect 3156 46752 3172 46816
rect 3236 46752 3252 46816
rect 3316 46752 3322 46816
rect 3006 46751 3322 46752
rect 8006 46816 8322 46817
rect 8006 46752 8012 46816
rect 8076 46752 8092 46816
rect 8156 46752 8172 46816
rect 8236 46752 8252 46816
rect 8316 46752 8322 46816
rect 8006 46751 8322 46752
rect 2346 46272 2662 46273
rect 2346 46208 2352 46272
rect 2416 46208 2432 46272
rect 2496 46208 2512 46272
rect 2576 46208 2592 46272
rect 2656 46208 2662 46272
rect 2346 46207 2662 46208
rect 7346 46272 7662 46273
rect 7346 46208 7352 46272
rect 7416 46208 7432 46272
rect 7496 46208 7512 46272
rect 7576 46208 7592 46272
rect 7656 46208 7662 46272
rect 7346 46207 7662 46208
rect 8385 46066 8451 46069
rect 9200 46066 10000 46096
rect 8385 46064 10000 46066
rect 8385 46008 8390 46064
rect 8446 46008 10000 46064
rect 8385 46006 10000 46008
rect 8385 46003 8451 46006
rect 9200 45976 10000 46006
rect 3006 45728 3322 45729
rect 3006 45664 3012 45728
rect 3076 45664 3092 45728
rect 3156 45664 3172 45728
rect 3236 45664 3252 45728
rect 3316 45664 3322 45728
rect 3006 45663 3322 45664
rect 8006 45728 8322 45729
rect 8006 45664 8012 45728
rect 8076 45664 8092 45728
rect 8156 45664 8172 45728
rect 8236 45664 8252 45728
rect 8316 45664 8322 45728
rect 8006 45663 8322 45664
rect 2346 45184 2662 45185
rect 2346 45120 2352 45184
rect 2416 45120 2432 45184
rect 2496 45120 2512 45184
rect 2576 45120 2592 45184
rect 2656 45120 2662 45184
rect 2346 45119 2662 45120
rect 7346 45184 7662 45185
rect 7346 45120 7352 45184
rect 7416 45120 7432 45184
rect 7496 45120 7512 45184
rect 7576 45120 7592 45184
rect 7656 45120 7662 45184
rect 7346 45119 7662 45120
rect 8385 44706 8451 44709
rect 9200 44706 10000 44736
rect 8385 44704 10000 44706
rect 8385 44648 8390 44704
rect 8446 44648 10000 44704
rect 8385 44646 10000 44648
rect 8385 44643 8451 44646
rect 3006 44640 3322 44641
rect 3006 44576 3012 44640
rect 3076 44576 3092 44640
rect 3156 44576 3172 44640
rect 3236 44576 3252 44640
rect 3316 44576 3322 44640
rect 3006 44575 3322 44576
rect 8006 44640 8322 44641
rect 8006 44576 8012 44640
rect 8076 44576 8092 44640
rect 8156 44576 8172 44640
rect 8236 44576 8252 44640
rect 8316 44576 8322 44640
rect 9200 44616 10000 44646
rect 8006 44575 8322 44576
rect 2346 44096 2662 44097
rect 2346 44032 2352 44096
rect 2416 44032 2432 44096
rect 2496 44032 2512 44096
rect 2576 44032 2592 44096
rect 2656 44032 2662 44096
rect 2346 44031 2662 44032
rect 7346 44096 7662 44097
rect 7346 44032 7352 44096
rect 7416 44032 7432 44096
rect 7496 44032 7512 44096
rect 7576 44032 7592 44096
rect 7656 44032 7662 44096
rect 7346 44031 7662 44032
rect 3006 43552 3322 43553
rect 3006 43488 3012 43552
rect 3076 43488 3092 43552
rect 3156 43488 3172 43552
rect 3236 43488 3252 43552
rect 3316 43488 3322 43552
rect 3006 43487 3322 43488
rect 8006 43552 8322 43553
rect 8006 43488 8012 43552
rect 8076 43488 8092 43552
rect 8156 43488 8172 43552
rect 8236 43488 8252 43552
rect 8316 43488 8322 43552
rect 8006 43487 8322 43488
rect 8845 43346 8911 43349
rect 9200 43346 10000 43376
rect 8845 43344 10000 43346
rect 8845 43288 8850 43344
rect 8906 43288 10000 43344
rect 8845 43286 10000 43288
rect 8845 43283 8911 43286
rect 9200 43256 10000 43286
rect 2346 43008 2662 43009
rect 2346 42944 2352 43008
rect 2416 42944 2432 43008
rect 2496 42944 2512 43008
rect 2576 42944 2592 43008
rect 2656 42944 2662 43008
rect 2346 42943 2662 42944
rect 7346 43008 7662 43009
rect 7346 42944 7352 43008
rect 7416 42944 7432 43008
rect 7496 42944 7512 43008
rect 7576 42944 7592 43008
rect 7656 42944 7662 43008
rect 7346 42943 7662 42944
rect 3006 42464 3322 42465
rect 3006 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3322 42464
rect 3006 42399 3322 42400
rect 8006 42464 8322 42465
rect 8006 42400 8012 42464
rect 8076 42400 8092 42464
rect 8156 42400 8172 42464
rect 8236 42400 8252 42464
rect 8316 42400 8322 42464
rect 8006 42399 8322 42400
rect 8385 41986 8451 41989
rect 9200 41986 10000 42016
rect 8385 41984 10000 41986
rect 8385 41928 8390 41984
rect 8446 41928 10000 41984
rect 8385 41926 10000 41928
rect 8385 41923 8451 41926
rect 2346 41920 2662 41921
rect 2346 41856 2352 41920
rect 2416 41856 2432 41920
rect 2496 41856 2512 41920
rect 2576 41856 2592 41920
rect 2656 41856 2662 41920
rect 2346 41855 2662 41856
rect 7346 41920 7662 41921
rect 7346 41856 7352 41920
rect 7416 41856 7432 41920
rect 7496 41856 7512 41920
rect 7576 41856 7592 41920
rect 7656 41856 7662 41920
rect 9200 41896 10000 41926
rect 7346 41855 7662 41856
rect 6177 41442 6243 41445
rect 6310 41442 6316 41444
rect 6177 41440 6316 41442
rect 6177 41384 6182 41440
rect 6238 41384 6316 41440
rect 6177 41382 6316 41384
rect 6177 41379 6243 41382
rect 6310 41380 6316 41382
rect 6380 41380 6386 41444
rect 3006 41376 3322 41377
rect 3006 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3322 41376
rect 3006 41311 3322 41312
rect 8006 41376 8322 41377
rect 8006 41312 8012 41376
rect 8076 41312 8092 41376
rect 8156 41312 8172 41376
rect 8236 41312 8252 41376
rect 8316 41312 8322 41376
rect 8006 41311 8322 41312
rect 2346 40832 2662 40833
rect 2346 40768 2352 40832
rect 2416 40768 2432 40832
rect 2496 40768 2512 40832
rect 2576 40768 2592 40832
rect 2656 40768 2662 40832
rect 2346 40767 2662 40768
rect 7346 40832 7662 40833
rect 7346 40768 7352 40832
rect 7416 40768 7432 40832
rect 7496 40768 7512 40832
rect 7576 40768 7592 40832
rect 7656 40768 7662 40832
rect 7346 40767 7662 40768
rect 8385 40626 8451 40629
rect 9200 40626 10000 40656
rect 8385 40624 10000 40626
rect 8385 40568 8390 40624
rect 8446 40568 10000 40624
rect 8385 40566 10000 40568
rect 8385 40563 8451 40566
rect 9200 40536 10000 40566
rect 3006 40288 3322 40289
rect 3006 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3322 40288
rect 3006 40223 3322 40224
rect 8006 40288 8322 40289
rect 8006 40224 8012 40288
rect 8076 40224 8092 40288
rect 8156 40224 8172 40288
rect 8236 40224 8252 40288
rect 8316 40224 8322 40288
rect 8006 40223 8322 40224
rect 5625 40082 5691 40085
rect 6678 40082 6684 40084
rect 5625 40080 6684 40082
rect 5625 40024 5630 40080
rect 5686 40024 6684 40080
rect 5625 40022 6684 40024
rect 5625 40019 5691 40022
rect 6678 40020 6684 40022
rect 6748 40020 6754 40084
rect 2346 39744 2662 39745
rect 2346 39680 2352 39744
rect 2416 39680 2432 39744
rect 2496 39680 2512 39744
rect 2576 39680 2592 39744
rect 2656 39680 2662 39744
rect 2346 39679 2662 39680
rect 7346 39744 7662 39745
rect 7346 39680 7352 39744
rect 7416 39680 7432 39744
rect 7496 39680 7512 39744
rect 7576 39680 7592 39744
rect 7656 39680 7662 39744
rect 7346 39679 7662 39680
rect 8385 39266 8451 39269
rect 9200 39266 10000 39296
rect 8385 39264 10000 39266
rect 8385 39208 8390 39264
rect 8446 39208 10000 39264
rect 8385 39206 10000 39208
rect 8385 39203 8451 39206
rect 3006 39200 3322 39201
rect 3006 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3322 39200
rect 3006 39135 3322 39136
rect 8006 39200 8322 39201
rect 8006 39136 8012 39200
rect 8076 39136 8092 39200
rect 8156 39136 8172 39200
rect 8236 39136 8252 39200
rect 8316 39136 8322 39200
rect 9200 39176 10000 39206
rect 8006 39135 8322 39136
rect 2346 38656 2662 38657
rect 2346 38592 2352 38656
rect 2416 38592 2432 38656
rect 2496 38592 2512 38656
rect 2576 38592 2592 38656
rect 2656 38592 2662 38656
rect 2346 38591 2662 38592
rect 7346 38656 7662 38657
rect 7346 38592 7352 38656
rect 7416 38592 7432 38656
rect 7496 38592 7512 38656
rect 7576 38592 7592 38656
rect 7656 38592 7662 38656
rect 7346 38591 7662 38592
rect 3006 38112 3322 38113
rect 3006 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3322 38112
rect 3006 38047 3322 38048
rect 8006 38112 8322 38113
rect 8006 38048 8012 38112
rect 8076 38048 8092 38112
rect 8156 38048 8172 38112
rect 8236 38048 8252 38112
rect 8316 38048 8322 38112
rect 8006 38047 8322 38048
rect 8385 37906 8451 37909
rect 9200 37906 10000 37936
rect 8385 37904 10000 37906
rect 8385 37848 8390 37904
rect 8446 37848 10000 37904
rect 8385 37846 10000 37848
rect 8385 37843 8451 37846
rect 9200 37816 10000 37846
rect 2346 37568 2662 37569
rect 2346 37504 2352 37568
rect 2416 37504 2432 37568
rect 2496 37504 2512 37568
rect 2576 37504 2592 37568
rect 2656 37504 2662 37568
rect 2346 37503 2662 37504
rect 7346 37568 7662 37569
rect 7346 37504 7352 37568
rect 7416 37504 7432 37568
rect 7496 37504 7512 37568
rect 7576 37504 7592 37568
rect 7656 37504 7662 37568
rect 7346 37503 7662 37504
rect 3006 37024 3322 37025
rect 3006 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3322 37024
rect 3006 36959 3322 36960
rect 8006 37024 8322 37025
rect 8006 36960 8012 37024
rect 8076 36960 8092 37024
rect 8156 36960 8172 37024
rect 8236 36960 8252 37024
rect 8316 36960 8322 37024
rect 8006 36959 8322 36960
rect 8385 36546 8451 36549
rect 9200 36546 10000 36576
rect 8385 36544 10000 36546
rect 8385 36488 8390 36544
rect 8446 36488 10000 36544
rect 8385 36486 10000 36488
rect 8385 36483 8451 36486
rect 2346 36480 2662 36481
rect 2346 36416 2352 36480
rect 2416 36416 2432 36480
rect 2496 36416 2512 36480
rect 2576 36416 2592 36480
rect 2656 36416 2662 36480
rect 2346 36415 2662 36416
rect 7346 36480 7662 36481
rect 7346 36416 7352 36480
rect 7416 36416 7432 36480
rect 7496 36416 7512 36480
rect 7576 36416 7592 36480
rect 7656 36416 7662 36480
rect 9200 36456 10000 36486
rect 7346 36415 7662 36416
rect 3006 35936 3322 35937
rect 3006 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3322 35936
rect 3006 35871 3322 35872
rect 8006 35936 8322 35937
rect 8006 35872 8012 35936
rect 8076 35872 8092 35936
rect 8156 35872 8172 35936
rect 8236 35872 8252 35936
rect 8316 35872 8322 35936
rect 8006 35871 8322 35872
rect 2346 35392 2662 35393
rect 2346 35328 2352 35392
rect 2416 35328 2432 35392
rect 2496 35328 2512 35392
rect 2576 35328 2592 35392
rect 2656 35328 2662 35392
rect 2346 35327 2662 35328
rect 7346 35392 7662 35393
rect 7346 35328 7352 35392
rect 7416 35328 7432 35392
rect 7496 35328 7512 35392
rect 7576 35328 7592 35392
rect 7656 35328 7662 35392
rect 7346 35327 7662 35328
rect 8385 35186 8451 35189
rect 9200 35186 10000 35216
rect 8385 35184 10000 35186
rect 8385 35128 8390 35184
rect 8446 35128 10000 35184
rect 8385 35126 10000 35128
rect 8385 35123 8451 35126
rect 9200 35096 10000 35126
rect 3006 34848 3322 34849
rect 3006 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3322 34848
rect 3006 34783 3322 34784
rect 8006 34848 8322 34849
rect 8006 34784 8012 34848
rect 8076 34784 8092 34848
rect 8156 34784 8172 34848
rect 8236 34784 8252 34848
rect 8316 34784 8322 34848
rect 8006 34783 8322 34784
rect 2346 34304 2662 34305
rect 2346 34240 2352 34304
rect 2416 34240 2432 34304
rect 2496 34240 2512 34304
rect 2576 34240 2592 34304
rect 2656 34240 2662 34304
rect 2346 34239 2662 34240
rect 7346 34304 7662 34305
rect 7346 34240 7352 34304
rect 7416 34240 7432 34304
rect 7496 34240 7512 34304
rect 7576 34240 7592 34304
rect 7656 34240 7662 34304
rect 7346 34239 7662 34240
rect 9200 33826 10000 33856
rect 8526 33766 10000 33826
rect 3006 33760 3322 33761
rect 3006 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3322 33760
rect 3006 33695 3322 33696
rect 8006 33760 8322 33761
rect 8006 33696 8012 33760
rect 8076 33696 8092 33760
rect 8156 33696 8172 33760
rect 8236 33696 8252 33760
rect 8316 33696 8322 33760
rect 8006 33695 8322 33696
rect 7741 33554 7807 33557
rect 8526 33554 8586 33766
rect 9200 33736 10000 33766
rect 7741 33552 8586 33554
rect 7741 33496 7746 33552
rect 7802 33496 8586 33552
rect 7741 33494 8586 33496
rect 7741 33491 7807 33494
rect 2346 33216 2662 33217
rect 2346 33152 2352 33216
rect 2416 33152 2432 33216
rect 2496 33152 2512 33216
rect 2576 33152 2592 33216
rect 2656 33152 2662 33216
rect 2346 33151 2662 33152
rect 7346 33216 7662 33217
rect 7346 33152 7352 33216
rect 7416 33152 7432 33216
rect 7496 33152 7512 33216
rect 7576 33152 7592 33216
rect 7656 33152 7662 33216
rect 7346 33151 7662 33152
rect 3006 32672 3322 32673
rect 3006 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3322 32672
rect 3006 32607 3322 32608
rect 8006 32672 8322 32673
rect 8006 32608 8012 32672
rect 8076 32608 8092 32672
rect 8156 32608 8172 32672
rect 8236 32608 8252 32672
rect 8316 32608 8322 32672
rect 8006 32607 8322 32608
rect 8661 32466 8727 32469
rect 9200 32466 10000 32496
rect 8661 32464 10000 32466
rect 8661 32408 8666 32464
rect 8722 32408 10000 32464
rect 8661 32406 10000 32408
rect 8661 32403 8727 32406
rect 9200 32376 10000 32406
rect 2346 32128 2662 32129
rect 2346 32064 2352 32128
rect 2416 32064 2432 32128
rect 2496 32064 2512 32128
rect 2576 32064 2592 32128
rect 2656 32064 2662 32128
rect 2346 32063 2662 32064
rect 7346 32128 7662 32129
rect 7346 32064 7352 32128
rect 7416 32064 7432 32128
rect 7496 32064 7512 32128
rect 7576 32064 7592 32128
rect 7656 32064 7662 32128
rect 7346 32063 7662 32064
rect 3006 31584 3322 31585
rect 3006 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3322 31584
rect 3006 31519 3322 31520
rect 8006 31584 8322 31585
rect 8006 31520 8012 31584
rect 8076 31520 8092 31584
rect 8156 31520 8172 31584
rect 8236 31520 8252 31584
rect 8316 31520 8322 31584
rect 8006 31519 8322 31520
rect 8385 31106 8451 31109
rect 9200 31106 10000 31136
rect 8385 31104 10000 31106
rect 8385 31048 8390 31104
rect 8446 31048 10000 31104
rect 8385 31046 10000 31048
rect 8385 31043 8451 31046
rect 2346 31040 2662 31041
rect 2346 30976 2352 31040
rect 2416 30976 2432 31040
rect 2496 30976 2512 31040
rect 2576 30976 2592 31040
rect 2656 30976 2662 31040
rect 2346 30975 2662 30976
rect 7346 31040 7662 31041
rect 7346 30976 7352 31040
rect 7416 30976 7432 31040
rect 7496 30976 7512 31040
rect 7576 30976 7592 31040
rect 7656 30976 7662 31040
rect 9200 31016 10000 31046
rect 7346 30975 7662 30976
rect 3006 30496 3322 30497
rect 3006 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3322 30496
rect 3006 30431 3322 30432
rect 8006 30496 8322 30497
rect 8006 30432 8012 30496
rect 8076 30432 8092 30496
rect 8156 30432 8172 30496
rect 8236 30432 8252 30496
rect 8316 30432 8322 30496
rect 8006 30431 8322 30432
rect 2346 29952 2662 29953
rect 2346 29888 2352 29952
rect 2416 29888 2432 29952
rect 2496 29888 2512 29952
rect 2576 29888 2592 29952
rect 2656 29888 2662 29952
rect 2346 29887 2662 29888
rect 7346 29952 7662 29953
rect 7346 29888 7352 29952
rect 7416 29888 7432 29952
rect 7496 29888 7512 29952
rect 7576 29888 7592 29952
rect 7656 29888 7662 29952
rect 7346 29887 7662 29888
rect 8385 29746 8451 29749
rect 9200 29746 10000 29776
rect 8385 29744 10000 29746
rect 8385 29688 8390 29744
rect 8446 29688 10000 29744
rect 8385 29686 10000 29688
rect 8385 29683 8451 29686
rect 9200 29656 10000 29686
rect 3006 29408 3322 29409
rect 3006 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3322 29408
rect 3006 29343 3322 29344
rect 8006 29408 8322 29409
rect 8006 29344 8012 29408
rect 8076 29344 8092 29408
rect 8156 29344 8172 29408
rect 8236 29344 8252 29408
rect 8316 29344 8322 29408
rect 8006 29343 8322 29344
rect 2346 28864 2662 28865
rect 2346 28800 2352 28864
rect 2416 28800 2432 28864
rect 2496 28800 2512 28864
rect 2576 28800 2592 28864
rect 2656 28800 2662 28864
rect 2346 28799 2662 28800
rect 7346 28864 7662 28865
rect 7346 28800 7352 28864
rect 7416 28800 7432 28864
rect 7496 28800 7512 28864
rect 7576 28800 7592 28864
rect 7656 28800 7662 28864
rect 7346 28799 7662 28800
rect 8385 28386 8451 28389
rect 9200 28386 10000 28416
rect 8385 28384 10000 28386
rect 8385 28328 8390 28384
rect 8446 28328 10000 28384
rect 8385 28326 10000 28328
rect 8385 28323 8451 28326
rect 3006 28320 3322 28321
rect 3006 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3322 28320
rect 3006 28255 3322 28256
rect 8006 28320 8322 28321
rect 8006 28256 8012 28320
rect 8076 28256 8092 28320
rect 8156 28256 8172 28320
rect 8236 28256 8252 28320
rect 8316 28256 8322 28320
rect 9200 28296 10000 28326
rect 8006 28255 8322 28256
rect 2346 27776 2662 27777
rect 2346 27712 2352 27776
rect 2416 27712 2432 27776
rect 2496 27712 2512 27776
rect 2576 27712 2592 27776
rect 2656 27712 2662 27776
rect 2346 27711 2662 27712
rect 7346 27776 7662 27777
rect 7346 27712 7352 27776
rect 7416 27712 7432 27776
rect 7496 27712 7512 27776
rect 7576 27712 7592 27776
rect 7656 27712 7662 27776
rect 7346 27711 7662 27712
rect 3006 27232 3322 27233
rect 3006 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3322 27232
rect 3006 27167 3322 27168
rect 8006 27232 8322 27233
rect 8006 27168 8012 27232
rect 8076 27168 8092 27232
rect 8156 27168 8172 27232
rect 8236 27168 8252 27232
rect 8316 27168 8322 27232
rect 8006 27167 8322 27168
rect 8845 27026 8911 27029
rect 9200 27026 10000 27056
rect 8845 27024 10000 27026
rect 8845 26968 8850 27024
rect 8906 26968 10000 27024
rect 8845 26966 10000 26968
rect 8845 26963 8911 26966
rect 9200 26936 10000 26966
rect 2346 26688 2662 26689
rect 2346 26624 2352 26688
rect 2416 26624 2432 26688
rect 2496 26624 2512 26688
rect 2576 26624 2592 26688
rect 2656 26624 2662 26688
rect 2346 26623 2662 26624
rect 7346 26688 7662 26689
rect 7346 26624 7352 26688
rect 7416 26624 7432 26688
rect 7496 26624 7512 26688
rect 7576 26624 7592 26688
rect 7656 26624 7662 26688
rect 7346 26623 7662 26624
rect 3006 26144 3322 26145
rect 3006 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3322 26144
rect 3006 26079 3322 26080
rect 8006 26144 8322 26145
rect 8006 26080 8012 26144
rect 8076 26080 8092 26144
rect 8156 26080 8172 26144
rect 8236 26080 8252 26144
rect 8316 26080 8322 26144
rect 8006 26079 8322 26080
rect 7741 25666 7807 25669
rect 9200 25666 10000 25696
rect 7741 25664 10000 25666
rect 7741 25608 7746 25664
rect 7802 25608 10000 25664
rect 7741 25606 10000 25608
rect 7741 25603 7807 25606
rect 2346 25600 2662 25601
rect 2346 25536 2352 25600
rect 2416 25536 2432 25600
rect 2496 25536 2512 25600
rect 2576 25536 2592 25600
rect 2656 25536 2662 25600
rect 2346 25535 2662 25536
rect 7346 25600 7662 25601
rect 7346 25536 7352 25600
rect 7416 25536 7432 25600
rect 7496 25536 7512 25600
rect 7576 25536 7592 25600
rect 7656 25536 7662 25600
rect 9200 25576 10000 25606
rect 7346 25535 7662 25536
rect 3006 25056 3322 25057
rect 3006 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3322 25056
rect 3006 24991 3322 24992
rect 8006 25056 8322 25057
rect 8006 24992 8012 25056
rect 8076 24992 8092 25056
rect 8156 24992 8172 25056
rect 8236 24992 8252 25056
rect 8316 24992 8322 25056
rect 8006 24991 8322 24992
rect 2346 24512 2662 24513
rect 2346 24448 2352 24512
rect 2416 24448 2432 24512
rect 2496 24448 2512 24512
rect 2576 24448 2592 24512
rect 2656 24448 2662 24512
rect 2346 24447 2662 24448
rect 7346 24512 7662 24513
rect 7346 24448 7352 24512
rect 7416 24448 7432 24512
rect 7496 24448 7512 24512
rect 7576 24448 7592 24512
rect 7656 24448 7662 24512
rect 7346 24447 7662 24448
rect 7373 24306 7439 24309
rect 9200 24306 10000 24336
rect 7373 24304 10000 24306
rect 7373 24248 7378 24304
rect 7434 24248 10000 24304
rect 7373 24246 10000 24248
rect 7373 24243 7439 24246
rect 9200 24216 10000 24246
rect 3006 23968 3322 23969
rect 3006 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3322 23968
rect 3006 23903 3322 23904
rect 8006 23968 8322 23969
rect 8006 23904 8012 23968
rect 8076 23904 8092 23968
rect 8156 23904 8172 23968
rect 8236 23904 8252 23968
rect 8316 23904 8322 23968
rect 8006 23903 8322 23904
rect 2346 23424 2662 23425
rect 2346 23360 2352 23424
rect 2416 23360 2432 23424
rect 2496 23360 2512 23424
rect 2576 23360 2592 23424
rect 2656 23360 2662 23424
rect 2346 23359 2662 23360
rect 7346 23424 7662 23425
rect 7346 23360 7352 23424
rect 7416 23360 7432 23424
rect 7496 23360 7512 23424
rect 7576 23360 7592 23424
rect 7656 23360 7662 23424
rect 7346 23359 7662 23360
rect 8385 22946 8451 22949
rect 9200 22946 10000 22976
rect 8385 22944 10000 22946
rect 8385 22888 8390 22944
rect 8446 22888 10000 22944
rect 8385 22886 10000 22888
rect 8385 22883 8451 22886
rect 3006 22880 3322 22881
rect 3006 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3322 22880
rect 3006 22815 3322 22816
rect 8006 22880 8322 22881
rect 8006 22816 8012 22880
rect 8076 22816 8092 22880
rect 8156 22816 8172 22880
rect 8236 22816 8252 22880
rect 8316 22816 8322 22880
rect 9200 22856 10000 22886
rect 8006 22815 8322 22816
rect 2346 22336 2662 22337
rect 2346 22272 2352 22336
rect 2416 22272 2432 22336
rect 2496 22272 2512 22336
rect 2576 22272 2592 22336
rect 2656 22272 2662 22336
rect 2346 22271 2662 22272
rect 7346 22336 7662 22337
rect 7346 22272 7352 22336
rect 7416 22272 7432 22336
rect 7496 22272 7512 22336
rect 7576 22272 7592 22336
rect 7656 22272 7662 22336
rect 7346 22271 7662 22272
rect 3006 21792 3322 21793
rect 3006 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3322 21792
rect 3006 21727 3322 21728
rect 8006 21792 8322 21793
rect 8006 21728 8012 21792
rect 8076 21728 8092 21792
rect 8156 21728 8172 21792
rect 8236 21728 8252 21792
rect 8316 21728 8322 21792
rect 8006 21727 8322 21728
rect 8293 21586 8359 21589
rect 9200 21586 10000 21616
rect 8293 21584 10000 21586
rect 8293 21528 8298 21584
rect 8354 21528 10000 21584
rect 8293 21526 10000 21528
rect 8293 21523 8359 21526
rect 9200 21496 10000 21526
rect 2346 21248 2662 21249
rect 2346 21184 2352 21248
rect 2416 21184 2432 21248
rect 2496 21184 2512 21248
rect 2576 21184 2592 21248
rect 2656 21184 2662 21248
rect 2346 21183 2662 21184
rect 7346 21248 7662 21249
rect 7346 21184 7352 21248
rect 7416 21184 7432 21248
rect 7496 21184 7512 21248
rect 7576 21184 7592 21248
rect 7656 21184 7662 21248
rect 7346 21183 7662 21184
rect 3006 20704 3322 20705
rect 3006 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3322 20704
rect 3006 20639 3322 20640
rect 8006 20704 8322 20705
rect 8006 20640 8012 20704
rect 8076 20640 8092 20704
rect 8156 20640 8172 20704
rect 8236 20640 8252 20704
rect 8316 20640 8322 20704
rect 8006 20639 8322 20640
rect 8293 20226 8359 20229
rect 9200 20226 10000 20256
rect 8293 20224 10000 20226
rect 8293 20168 8298 20224
rect 8354 20168 10000 20224
rect 8293 20166 10000 20168
rect 8293 20163 8359 20166
rect 2346 20160 2662 20161
rect 2346 20096 2352 20160
rect 2416 20096 2432 20160
rect 2496 20096 2512 20160
rect 2576 20096 2592 20160
rect 2656 20096 2662 20160
rect 2346 20095 2662 20096
rect 7346 20160 7662 20161
rect 7346 20096 7352 20160
rect 7416 20096 7432 20160
rect 7496 20096 7512 20160
rect 7576 20096 7592 20160
rect 7656 20096 7662 20160
rect 9200 20136 10000 20166
rect 7346 20095 7662 20096
rect 3006 19616 3322 19617
rect 3006 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3322 19616
rect 3006 19551 3322 19552
rect 8006 19616 8322 19617
rect 8006 19552 8012 19616
rect 8076 19552 8092 19616
rect 8156 19552 8172 19616
rect 8236 19552 8252 19616
rect 8316 19552 8322 19616
rect 8006 19551 8322 19552
rect 2346 19072 2662 19073
rect 2346 19008 2352 19072
rect 2416 19008 2432 19072
rect 2496 19008 2512 19072
rect 2576 19008 2592 19072
rect 2656 19008 2662 19072
rect 2346 19007 2662 19008
rect 7346 19072 7662 19073
rect 7346 19008 7352 19072
rect 7416 19008 7432 19072
rect 7496 19008 7512 19072
rect 7576 19008 7592 19072
rect 7656 19008 7662 19072
rect 7346 19007 7662 19008
rect 8201 18866 8267 18869
rect 9200 18866 10000 18896
rect 8201 18864 10000 18866
rect 8201 18808 8206 18864
rect 8262 18808 10000 18864
rect 8201 18806 10000 18808
rect 8201 18803 8267 18806
rect 9200 18776 10000 18806
rect 3006 18528 3322 18529
rect 3006 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3322 18528
rect 3006 18463 3322 18464
rect 8006 18528 8322 18529
rect 8006 18464 8012 18528
rect 8076 18464 8092 18528
rect 8156 18464 8172 18528
rect 8236 18464 8252 18528
rect 8316 18464 8322 18528
rect 8006 18463 8322 18464
rect 2346 17984 2662 17985
rect 2346 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2662 17984
rect 2346 17919 2662 17920
rect 7346 17984 7662 17985
rect 7346 17920 7352 17984
rect 7416 17920 7432 17984
rect 7496 17920 7512 17984
rect 7576 17920 7592 17984
rect 7656 17920 7662 17984
rect 7346 17919 7662 17920
rect 8477 17506 8543 17509
rect 9200 17506 10000 17536
rect 8477 17504 10000 17506
rect 8477 17448 8482 17504
rect 8538 17448 10000 17504
rect 8477 17446 10000 17448
rect 8477 17443 8543 17446
rect 3006 17440 3322 17441
rect 3006 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3322 17440
rect 3006 17375 3322 17376
rect 8006 17440 8322 17441
rect 8006 17376 8012 17440
rect 8076 17376 8092 17440
rect 8156 17376 8172 17440
rect 8236 17376 8252 17440
rect 8316 17376 8322 17440
rect 9200 17416 10000 17446
rect 8006 17375 8322 17376
rect 2346 16896 2662 16897
rect 2346 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2662 16896
rect 2346 16831 2662 16832
rect 7346 16896 7662 16897
rect 7346 16832 7352 16896
rect 7416 16832 7432 16896
rect 7496 16832 7512 16896
rect 7576 16832 7592 16896
rect 7656 16832 7662 16896
rect 7346 16831 7662 16832
rect 3006 16352 3322 16353
rect 3006 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3322 16352
rect 3006 16287 3322 16288
rect 8006 16352 8322 16353
rect 8006 16288 8012 16352
rect 8076 16288 8092 16352
rect 8156 16288 8172 16352
rect 8236 16288 8252 16352
rect 8316 16288 8322 16352
rect 8006 16287 8322 16288
rect 6729 16146 6795 16149
rect 9200 16146 10000 16176
rect 6729 16144 10000 16146
rect 6729 16088 6734 16144
rect 6790 16088 10000 16144
rect 6729 16086 10000 16088
rect 6729 16083 6795 16086
rect 9200 16056 10000 16086
rect 2346 15808 2662 15809
rect 2346 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2662 15808
rect 2346 15743 2662 15744
rect 7346 15808 7662 15809
rect 7346 15744 7352 15808
rect 7416 15744 7432 15808
rect 7496 15744 7512 15808
rect 7576 15744 7592 15808
rect 7656 15744 7662 15808
rect 7346 15743 7662 15744
rect 3006 15264 3322 15265
rect 3006 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3322 15264
rect 3006 15199 3322 15200
rect 8006 15264 8322 15265
rect 8006 15200 8012 15264
rect 8076 15200 8092 15264
rect 8156 15200 8172 15264
rect 8236 15200 8252 15264
rect 8316 15200 8322 15264
rect 8006 15199 8322 15200
rect 8845 14786 8911 14789
rect 9200 14786 10000 14816
rect 8845 14784 10000 14786
rect 8845 14728 8850 14784
rect 8906 14728 10000 14784
rect 8845 14726 10000 14728
rect 8845 14723 8911 14726
rect 2346 14720 2662 14721
rect 2346 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2662 14720
rect 2346 14655 2662 14656
rect 7346 14720 7662 14721
rect 7346 14656 7352 14720
rect 7416 14656 7432 14720
rect 7496 14656 7512 14720
rect 7576 14656 7592 14720
rect 7656 14656 7662 14720
rect 9200 14696 10000 14726
rect 7346 14655 7662 14656
rect 3006 14176 3322 14177
rect 3006 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3322 14176
rect 3006 14111 3322 14112
rect 8006 14176 8322 14177
rect 8006 14112 8012 14176
rect 8076 14112 8092 14176
rect 8156 14112 8172 14176
rect 8236 14112 8252 14176
rect 8316 14112 8322 14176
rect 8006 14111 8322 14112
rect 2346 13632 2662 13633
rect 2346 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2662 13632
rect 2346 13567 2662 13568
rect 7346 13632 7662 13633
rect 7346 13568 7352 13632
rect 7416 13568 7432 13632
rect 7496 13568 7512 13632
rect 7576 13568 7592 13632
rect 7656 13568 7662 13632
rect 7346 13567 7662 13568
rect 8293 13426 8359 13429
rect 9200 13426 10000 13456
rect 8293 13424 10000 13426
rect 8293 13368 8298 13424
rect 8354 13368 10000 13424
rect 8293 13366 10000 13368
rect 8293 13363 8359 13366
rect 9200 13336 10000 13366
rect 3006 13088 3322 13089
rect 3006 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3322 13088
rect 3006 13023 3322 13024
rect 8006 13088 8322 13089
rect 8006 13024 8012 13088
rect 8076 13024 8092 13088
rect 8156 13024 8172 13088
rect 8236 13024 8252 13088
rect 8316 13024 8322 13088
rect 8006 13023 8322 13024
rect 2346 12544 2662 12545
rect 2346 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2662 12544
rect 2346 12479 2662 12480
rect 7346 12544 7662 12545
rect 7346 12480 7352 12544
rect 7416 12480 7432 12544
rect 7496 12480 7512 12544
rect 7576 12480 7592 12544
rect 7656 12480 7662 12544
rect 7346 12479 7662 12480
rect 8477 12066 8543 12069
rect 9200 12066 10000 12096
rect 8477 12064 10000 12066
rect 8477 12008 8482 12064
rect 8538 12008 10000 12064
rect 8477 12006 10000 12008
rect 8477 12003 8543 12006
rect 3006 12000 3322 12001
rect 3006 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3322 12000
rect 3006 11935 3322 11936
rect 8006 12000 8322 12001
rect 8006 11936 8012 12000
rect 8076 11936 8092 12000
rect 8156 11936 8172 12000
rect 8236 11936 8252 12000
rect 8316 11936 8322 12000
rect 9200 11976 10000 12006
rect 8006 11935 8322 11936
rect 2346 11456 2662 11457
rect 2346 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2662 11456
rect 2346 11391 2662 11392
rect 7346 11456 7662 11457
rect 7346 11392 7352 11456
rect 7416 11392 7432 11456
rect 7496 11392 7512 11456
rect 7576 11392 7592 11456
rect 7656 11392 7662 11456
rect 7346 11391 7662 11392
rect 3006 10912 3322 10913
rect 3006 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3322 10912
rect 3006 10847 3322 10848
rect 8006 10912 8322 10913
rect 8006 10848 8012 10912
rect 8076 10848 8092 10912
rect 8156 10848 8172 10912
rect 8236 10848 8252 10912
rect 8316 10848 8322 10912
rect 8006 10847 8322 10848
rect 7925 10706 7991 10709
rect 9200 10706 10000 10736
rect 7925 10704 10000 10706
rect 7925 10648 7930 10704
rect 7986 10648 10000 10704
rect 7925 10646 10000 10648
rect 7925 10643 7991 10646
rect 9200 10616 10000 10646
rect 2346 10368 2662 10369
rect 2346 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2662 10368
rect 2346 10303 2662 10304
rect 7346 10368 7662 10369
rect 7346 10304 7352 10368
rect 7416 10304 7432 10368
rect 7496 10304 7512 10368
rect 7576 10304 7592 10368
rect 7656 10304 7662 10368
rect 7346 10303 7662 10304
rect 3006 9824 3322 9825
rect 3006 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3322 9824
rect 3006 9759 3322 9760
rect 8006 9824 8322 9825
rect 8006 9760 8012 9824
rect 8076 9760 8092 9824
rect 8156 9760 8172 9824
rect 8236 9760 8252 9824
rect 8316 9760 8322 9824
rect 8006 9759 8322 9760
rect 8293 9346 8359 9349
rect 9200 9346 10000 9376
rect 8293 9344 10000 9346
rect 8293 9288 8298 9344
rect 8354 9288 10000 9344
rect 8293 9286 10000 9288
rect 8293 9283 8359 9286
rect 2346 9280 2662 9281
rect 2346 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2662 9280
rect 2346 9215 2662 9216
rect 7346 9280 7662 9281
rect 7346 9216 7352 9280
rect 7416 9216 7432 9280
rect 7496 9216 7512 9280
rect 7576 9216 7592 9280
rect 7656 9216 7662 9280
rect 9200 9256 10000 9286
rect 7346 9215 7662 9216
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 8006 8736 8322 8737
rect 8006 8672 8012 8736
rect 8076 8672 8092 8736
rect 8156 8672 8172 8736
rect 8236 8672 8252 8736
rect 8316 8672 8322 8736
rect 8006 8671 8322 8672
rect 2346 8192 2662 8193
rect 2346 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2662 8192
rect 2346 8127 2662 8128
rect 7346 8192 7662 8193
rect 7346 8128 7352 8192
rect 7416 8128 7432 8192
rect 7496 8128 7512 8192
rect 7576 8128 7592 8192
rect 7656 8128 7662 8192
rect 7346 8127 7662 8128
rect 7005 7986 7071 7989
rect 9200 7986 10000 8016
rect 7005 7984 10000 7986
rect 7005 7928 7010 7984
rect 7066 7928 10000 7984
rect 7005 7926 10000 7928
rect 7005 7923 7071 7926
rect 9200 7896 10000 7926
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 8006 7648 8322 7649
rect 8006 7584 8012 7648
rect 8076 7584 8092 7648
rect 8156 7584 8172 7648
rect 8236 7584 8252 7648
rect 8316 7584 8322 7648
rect 8006 7583 8322 7584
rect 2346 7104 2662 7105
rect 2346 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2662 7104
rect 2346 7039 2662 7040
rect 7346 7104 7662 7105
rect 7346 7040 7352 7104
rect 7416 7040 7432 7104
rect 7496 7040 7512 7104
rect 7576 7040 7592 7104
rect 7656 7040 7662 7104
rect 7346 7039 7662 7040
rect 6310 6836 6316 6900
rect 6380 6898 6386 6900
rect 7649 6898 7715 6901
rect 6380 6896 7715 6898
rect 6380 6840 7654 6896
rect 7710 6840 7715 6896
rect 6380 6838 7715 6840
rect 6380 6836 6386 6838
rect 7649 6835 7715 6838
rect 8845 6626 8911 6629
rect 9200 6626 10000 6656
rect 8845 6624 10000 6626
rect 8845 6568 8850 6624
rect 8906 6568 10000 6624
rect 8845 6566 10000 6568
rect 8845 6563 8911 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 8006 6560 8322 6561
rect 8006 6496 8012 6560
rect 8076 6496 8092 6560
rect 8156 6496 8172 6560
rect 8236 6496 8252 6560
rect 8316 6496 8322 6560
rect 9200 6536 10000 6566
rect 8006 6495 8322 6496
rect 2346 6016 2662 6017
rect 2346 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2662 6016
rect 2346 5951 2662 5952
rect 7346 6016 7662 6017
rect 7346 5952 7352 6016
rect 7416 5952 7432 6016
rect 7496 5952 7512 6016
rect 7576 5952 7592 6016
rect 7656 5952 7662 6016
rect 7346 5951 7662 5952
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 8006 5472 8322 5473
rect 8006 5408 8012 5472
rect 8076 5408 8092 5472
rect 8156 5408 8172 5472
rect 8236 5408 8252 5472
rect 8316 5408 8322 5472
rect 8006 5407 8322 5408
rect 2346 4928 2662 4929
rect 2346 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2662 4928
rect 2346 4863 2662 4864
rect 7346 4928 7662 4929
rect 7346 4864 7352 4928
rect 7416 4864 7432 4928
rect 7496 4864 7512 4928
rect 7576 4864 7592 4928
rect 7656 4864 7662 4928
rect 7346 4863 7662 4864
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 8006 4384 8322 4385
rect 8006 4320 8012 4384
rect 8076 4320 8092 4384
rect 8156 4320 8172 4384
rect 8236 4320 8252 4384
rect 8316 4320 8322 4384
rect 8006 4319 8322 4320
rect 2346 3840 2662 3841
rect 2346 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2662 3840
rect 2346 3775 2662 3776
rect 7346 3840 7662 3841
rect 7346 3776 7352 3840
rect 7416 3776 7432 3840
rect 7496 3776 7512 3840
rect 7576 3776 7592 3840
rect 7656 3776 7662 3840
rect 7346 3775 7662 3776
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 8006 3296 8322 3297
rect 8006 3232 8012 3296
rect 8076 3232 8092 3296
rect 8156 3232 8172 3296
rect 8236 3232 8252 3296
rect 8316 3232 8322 3296
rect 8006 3231 8322 3232
rect 2346 2752 2662 2753
rect 2346 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2662 2752
rect 2346 2687 2662 2688
rect 7346 2752 7662 2753
rect 7346 2688 7352 2752
rect 7416 2688 7432 2752
rect 7496 2688 7512 2752
rect 7576 2688 7592 2752
rect 7656 2688 7662 2752
rect 7346 2687 7662 2688
rect 6637 2684 6703 2685
rect 6637 2680 6684 2684
rect 6748 2682 6754 2684
rect 6637 2624 6642 2680
rect 6637 2620 6684 2624
rect 6748 2622 6794 2682
rect 6748 2620 6754 2622
rect 6637 2619 6703 2620
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 8006 2208 8322 2209
rect 8006 2144 8012 2208
rect 8076 2144 8092 2208
rect 8156 2144 8172 2208
rect 8236 2144 8252 2208
rect 8316 2144 8322 2208
rect 8006 2143 8322 2144
<< via3 >>
rect 2352 77820 2416 77824
rect 2352 77764 2356 77820
rect 2356 77764 2412 77820
rect 2412 77764 2416 77820
rect 2352 77760 2416 77764
rect 2432 77820 2496 77824
rect 2432 77764 2436 77820
rect 2436 77764 2492 77820
rect 2492 77764 2496 77820
rect 2432 77760 2496 77764
rect 2512 77820 2576 77824
rect 2512 77764 2516 77820
rect 2516 77764 2572 77820
rect 2572 77764 2576 77820
rect 2512 77760 2576 77764
rect 2592 77820 2656 77824
rect 2592 77764 2596 77820
rect 2596 77764 2652 77820
rect 2652 77764 2656 77820
rect 2592 77760 2656 77764
rect 7352 77820 7416 77824
rect 7352 77764 7356 77820
rect 7356 77764 7412 77820
rect 7412 77764 7416 77820
rect 7352 77760 7416 77764
rect 7432 77820 7496 77824
rect 7432 77764 7436 77820
rect 7436 77764 7492 77820
rect 7492 77764 7496 77820
rect 7432 77760 7496 77764
rect 7512 77820 7576 77824
rect 7512 77764 7516 77820
rect 7516 77764 7572 77820
rect 7572 77764 7576 77820
rect 7512 77760 7576 77764
rect 7592 77820 7656 77824
rect 7592 77764 7596 77820
rect 7596 77764 7652 77820
rect 7652 77764 7656 77820
rect 7592 77760 7656 77764
rect 3012 77276 3076 77280
rect 3012 77220 3016 77276
rect 3016 77220 3072 77276
rect 3072 77220 3076 77276
rect 3012 77216 3076 77220
rect 3092 77276 3156 77280
rect 3092 77220 3096 77276
rect 3096 77220 3152 77276
rect 3152 77220 3156 77276
rect 3092 77216 3156 77220
rect 3172 77276 3236 77280
rect 3172 77220 3176 77276
rect 3176 77220 3232 77276
rect 3232 77220 3236 77276
rect 3172 77216 3236 77220
rect 3252 77276 3316 77280
rect 3252 77220 3256 77276
rect 3256 77220 3312 77276
rect 3312 77220 3316 77276
rect 3252 77216 3316 77220
rect 8012 77276 8076 77280
rect 8012 77220 8016 77276
rect 8016 77220 8072 77276
rect 8072 77220 8076 77276
rect 8012 77216 8076 77220
rect 8092 77276 8156 77280
rect 8092 77220 8096 77276
rect 8096 77220 8152 77276
rect 8152 77220 8156 77276
rect 8092 77216 8156 77220
rect 8172 77276 8236 77280
rect 8172 77220 8176 77276
rect 8176 77220 8232 77276
rect 8232 77220 8236 77276
rect 8172 77216 8236 77220
rect 8252 77276 8316 77280
rect 8252 77220 8256 77276
rect 8256 77220 8312 77276
rect 8312 77220 8316 77276
rect 8252 77216 8316 77220
rect 2352 76732 2416 76736
rect 2352 76676 2356 76732
rect 2356 76676 2412 76732
rect 2412 76676 2416 76732
rect 2352 76672 2416 76676
rect 2432 76732 2496 76736
rect 2432 76676 2436 76732
rect 2436 76676 2492 76732
rect 2492 76676 2496 76732
rect 2432 76672 2496 76676
rect 2512 76732 2576 76736
rect 2512 76676 2516 76732
rect 2516 76676 2572 76732
rect 2572 76676 2576 76732
rect 2512 76672 2576 76676
rect 2592 76732 2656 76736
rect 2592 76676 2596 76732
rect 2596 76676 2652 76732
rect 2652 76676 2656 76732
rect 2592 76672 2656 76676
rect 7352 76732 7416 76736
rect 7352 76676 7356 76732
rect 7356 76676 7412 76732
rect 7412 76676 7416 76732
rect 7352 76672 7416 76676
rect 7432 76732 7496 76736
rect 7432 76676 7436 76732
rect 7436 76676 7492 76732
rect 7492 76676 7496 76732
rect 7432 76672 7496 76676
rect 7512 76732 7576 76736
rect 7512 76676 7516 76732
rect 7516 76676 7572 76732
rect 7572 76676 7576 76732
rect 7512 76672 7576 76676
rect 7592 76732 7656 76736
rect 7592 76676 7596 76732
rect 7596 76676 7652 76732
rect 7652 76676 7656 76732
rect 7592 76672 7656 76676
rect 3012 76188 3076 76192
rect 3012 76132 3016 76188
rect 3016 76132 3072 76188
rect 3072 76132 3076 76188
rect 3012 76128 3076 76132
rect 3092 76188 3156 76192
rect 3092 76132 3096 76188
rect 3096 76132 3152 76188
rect 3152 76132 3156 76188
rect 3092 76128 3156 76132
rect 3172 76188 3236 76192
rect 3172 76132 3176 76188
rect 3176 76132 3232 76188
rect 3232 76132 3236 76188
rect 3172 76128 3236 76132
rect 3252 76188 3316 76192
rect 3252 76132 3256 76188
rect 3256 76132 3312 76188
rect 3312 76132 3316 76188
rect 3252 76128 3316 76132
rect 8012 76188 8076 76192
rect 8012 76132 8016 76188
rect 8016 76132 8072 76188
rect 8072 76132 8076 76188
rect 8012 76128 8076 76132
rect 8092 76188 8156 76192
rect 8092 76132 8096 76188
rect 8096 76132 8152 76188
rect 8152 76132 8156 76188
rect 8092 76128 8156 76132
rect 8172 76188 8236 76192
rect 8172 76132 8176 76188
rect 8176 76132 8232 76188
rect 8232 76132 8236 76188
rect 8172 76128 8236 76132
rect 8252 76188 8316 76192
rect 8252 76132 8256 76188
rect 8256 76132 8312 76188
rect 8312 76132 8316 76188
rect 8252 76128 8316 76132
rect 2352 75644 2416 75648
rect 2352 75588 2356 75644
rect 2356 75588 2412 75644
rect 2412 75588 2416 75644
rect 2352 75584 2416 75588
rect 2432 75644 2496 75648
rect 2432 75588 2436 75644
rect 2436 75588 2492 75644
rect 2492 75588 2496 75644
rect 2432 75584 2496 75588
rect 2512 75644 2576 75648
rect 2512 75588 2516 75644
rect 2516 75588 2572 75644
rect 2572 75588 2576 75644
rect 2512 75584 2576 75588
rect 2592 75644 2656 75648
rect 2592 75588 2596 75644
rect 2596 75588 2652 75644
rect 2652 75588 2656 75644
rect 2592 75584 2656 75588
rect 7352 75644 7416 75648
rect 7352 75588 7356 75644
rect 7356 75588 7412 75644
rect 7412 75588 7416 75644
rect 7352 75584 7416 75588
rect 7432 75644 7496 75648
rect 7432 75588 7436 75644
rect 7436 75588 7492 75644
rect 7492 75588 7496 75644
rect 7432 75584 7496 75588
rect 7512 75644 7576 75648
rect 7512 75588 7516 75644
rect 7516 75588 7572 75644
rect 7572 75588 7576 75644
rect 7512 75584 7576 75588
rect 7592 75644 7656 75648
rect 7592 75588 7596 75644
rect 7596 75588 7652 75644
rect 7652 75588 7656 75644
rect 7592 75584 7656 75588
rect 3012 75100 3076 75104
rect 3012 75044 3016 75100
rect 3016 75044 3072 75100
rect 3072 75044 3076 75100
rect 3012 75040 3076 75044
rect 3092 75100 3156 75104
rect 3092 75044 3096 75100
rect 3096 75044 3152 75100
rect 3152 75044 3156 75100
rect 3092 75040 3156 75044
rect 3172 75100 3236 75104
rect 3172 75044 3176 75100
rect 3176 75044 3232 75100
rect 3232 75044 3236 75100
rect 3172 75040 3236 75044
rect 3252 75100 3316 75104
rect 3252 75044 3256 75100
rect 3256 75044 3312 75100
rect 3312 75044 3316 75100
rect 3252 75040 3316 75044
rect 8012 75100 8076 75104
rect 8012 75044 8016 75100
rect 8016 75044 8072 75100
rect 8072 75044 8076 75100
rect 8012 75040 8076 75044
rect 8092 75100 8156 75104
rect 8092 75044 8096 75100
rect 8096 75044 8152 75100
rect 8152 75044 8156 75100
rect 8092 75040 8156 75044
rect 8172 75100 8236 75104
rect 8172 75044 8176 75100
rect 8176 75044 8232 75100
rect 8232 75044 8236 75100
rect 8172 75040 8236 75044
rect 8252 75100 8316 75104
rect 8252 75044 8256 75100
rect 8256 75044 8312 75100
rect 8312 75044 8316 75100
rect 8252 75040 8316 75044
rect 2352 74556 2416 74560
rect 2352 74500 2356 74556
rect 2356 74500 2412 74556
rect 2412 74500 2416 74556
rect 2352 74496 2416 74500
rect 2432 74556 2496 74560
rect 2432 74500 2436 74556
rect 2436 74500 2492 74556
rect 2492 74500 2496 74556
rect 2432 74496 2496 74500
rect 2512 74556 2576 74560
rect 2512 74500 2516 74556
rect 2516 74500 2572 74556
rect 2572 74500 2576 74556
rect 2512 74496 2576 74500
rect 2592 74556 2656 74560
rect 2592 74500 2596 74556
rect 2596 74500 2652 74556
rect 2652 74500 2656 74556
rect 2592 74496 2656 74500
rect 7352 74556 7416 74560
rect 7352 74500 7356 74556
rect 7356 74500 7412 74556
rect 7412 74500 7416 74556
rect 7352 74496 7416 74500
rect 7432 74556 7496 74560
rect 7432 74500 7436 74556
rect 7436 74500 7492 74556
rect 7492 74500 7496 74556
rect 7432 74496 7496 74500
rect 7512 74556 7576 74560
rect 7512 74500 7516 74556
rect 7516 74500 7572 74556
rect 7572 74500 7576 74556
rect 7512 74496 7576 74500
rect 7592 74556 7656 74560
rect 7592 74500 7596 74556
rect 7596 74500 7652 74556
rect 7652 74500 7656 74556
rect 7592 74496 7656 74500
rect 3012 74012 3076 74016
rect 3012 73956 3016 74012
rect 3016 73956 3072 74012
rect 3072 73956 3076 74012
rect 3012 73952 3076 73956
rect 3092 74012 3156 74016
rect 3092 73956 3096 74012
rect 3096 73956 3152 74012
rect 3152 73956 3156 74012
rect 3092 73952 3156 73956
rect 3172 74012 3236 74016
rect 3172 73956 3176 74012
rect 3176 73956 3232 74012
rect 3232 73956 3236 74012
rect 3172 73952 3236 73956
rect 3252 74012 3316 74016
rect 3252 73956 3256 74012
rect 3256 73956 3312 74012
rect 3312 73956 3316 74012
rect 3252 73952 3316 73956
rect 8012 74012 8076 74016
rect 8012 73956 8016 74012
rect 8016 73956 8072 74012
rect 8072 73956 8076 74012
rect 8012 73952 8076 73956
rect 8092 74012 8156 74016
rect 8092 73956 8096 74012
rect 8096 73956 8152 74012
rect 8152 73956 8156 74012
rect 8092 73952 8156 73956
rect 8172 74012 8236 74016
rect 8172 73956 8176 74012
rect 8176 73956 8232 74012
rect 8232 73956 8236 74012
rect 8172 73952 8236 73956
rect 8252 74012 8316 74016
rect 8252 73956 8256 74012
rect 8256 73956 8312 74012
rect 8312 73956 8316 74012
rect 8252 73952 8316 73956
rect 2352 73468 2416 73472
rect 2352 73412 2356 73468
rect 2356 73412 2412 73468
rect 2412 73412 2416 73468
rect 2352 73408 2416 73412
rect 2432 73468 2496 73472
rect 2432 73412 2436 73468
rect 2436 73412 2492 73468
rect 2492 73412 2496 73468
rect 2432 73408 2496 73412
rect 2512 73468 2576 73472
rect 2512 73412 2516 73468
rect 2516 73412 2572 73468
rect 2572 73412 2576 73468
rect 2512 73408 2576 73412
rect 2592 73468 2656 73472
rect 2592 73412 2596 73468
rect 2596 73412 2652 73468
rect 2652 73412 2656 73468
rect 2592 73408 2656 73412
rect 7352 73468 7416 73472
rect 7352 73412 7356 73468
rect 7356 73412 7412 73468
rect 7412 73412 7416 73468
rect 7352 73408 7416 73412
rect 7432 73468 7496 73472
rect 7432 73412 7436 73468
rect 7436 73412 7492 73468
rect 7492 73412 7496 73468
rect 7432 73408 7496 73412
rect 7512 73468 7576 73472
rect 7512 73412 7516 73468
rect 7516 73412 7572 73468
rect 7572 73412 7576 73468
rect 7512 73408 7576 73412
rect 7592 73468 7656 73472
rect 7592 73412 7596 73468
rect 7596 73412 7652 73468
rect 7652 73412 7656 73468
rect 7592 73408 7656 73412
rect 3012 72924 3076 72928
rect 3012 72868 3016 72924
rect 3016 72868 3072 72924
rect 3072 72868 3076 72924
rect 3012 72864 3076 72868
rect 3092 72924 3156 72928
rect 3092 72868 3096 72924
rect 3096 72868 3152 72924
rect 3152 72868 3156 72924
rect 3092 72864 3156 72868
rect 3172 72924 3236 72928
rect 3172 72868 3176 72924
rect 3176 72868 3232 72924
rect 3232 72868 3236 72924
rect 3172 72864 3236 72868
rect 3252 72924 3316 72928
rect 3252 72868 3256 72924
rect 3256 72868 3312 72924
rect 3312 72868 3316 72924
rect 3252 72864 3316 72868
rect 8012 72924 8076 72928
rect 8012 72868 8016 72924
rect 8016 72868 8072 72924
rect 8072 72868 8076 72924
rect 8012 72864 8076 72868
rect 8092 72924 8156 72928
rect 8092 72868 8096 72924
rect 8096 72868 8152 72924
rect 8152 72868 8156 72924
rect 8092 72864 8156 72868
rect 8172 72924 8236 72928
rect 8172 72868 8176 72924
rect 8176 72868 8232 72924
rect 8232 72868 8236 72924
rect 8172 72864 8236 72868
rect 8252 72924 8316 72928
rect 8252 72868 8256 72924
rect 8256 72868 8312 72924
rect 8312 72868 8316 72924
rect 8252 72864 8316 72868
rect 2352 72380 2416 72384
rect 2352 72324 2356 72380
rect 2356 72324 2412 72380
rect 2412 72324 2416 72380
rect 2352 72320 2416 72324
rect 2432 72380 2496 72384
rect 2432 72324 2436 72380
rect 2436 72324 2492 72380
rect 2492 72324 2496 72380
rect 2432 72320 2496 72324
rect 2512 72380 2576 72384
rect 2512 72324 2516 72380
rect 2516 72324 2572 72380
rect 2572 72324 2576 72380
rect 2512 72320 2576 72324
rect 2592 72380 2656 72384
rect 2592 72324 2596 72380
rect 2596 72324 2652 72380
rect 2652 72324 2656 72380
rect 2592 72320 2656 72324
rect 7352 72380 7416 72384
rect 7352 72324 7356 72380
rect 7356 72324 7412 72380
rect 7412 72324 7416 72380
rect 7352 72320 7416 72324
rect 7432 72380 7496 72384
rect 7432 72324 7436 72380
rect 7436 72324 7492 72380
rect 7492 72324 7496 72380
rect 7432 72320 7496 72324
rect 7512 72380 7576 72384
rect 7512 72324 7516 72380
rect 7516 72324 7572 72380
rect 7572 72324 7576 72380
rect 7512 72320 7576 72324
rect 7592 72380 7656 72384
rect 7592 72324 7596 72380
rect 7596 72324 7652 72380
rect 7652 72324 7656 72380
rect 7592 72320 7656 72324
rect 3012 71836 3076 71840
rect 3012 71780 3016 71836
rect 3016 71780 3072 71836
rect 3072 71780 3076 71836
rect 3012 71776 3076 71780
rect 3092 71836 3156 71840
rect 3092 71780 3096 71836
rect 3096 71780 3152 71836
rect 3152 71780 3156 71836
rect 3092 71776 3156 71780
rect 3172 71836 3236 71840
rect 3172 71780 3176 71836
rect 3176 71780 3232 71836
rect 3232 71780 3236 71836
rect 3172 71776 3236 71780
rect 3252 71836 3316 71840
rect 3252 71780 3256 71836
rect 3256 71780 3312 71836
rect 3312 71780 3316 71836
rect 3252 71776 3316 71780
rect 8012 71836 8076 71840
rect 8012 71780 8016 71836
rect 8016 71780 8072 71836
rect 8072 71780 8076 71836
rect 8012 71776 8076 71780
rect 8092 71836 8156 71840
rect 8092 71780 8096 71836
rect 8096 71780 8152 71836
rect 8152 71780 8156 71836
rect 8092 71776 8156 71780
rect 8172 71836 8236 71840
rect 8172 71780 8176 71836
rect 8176 71780 8232 71836
rect 8232 71780 8236 71836
rect 8172 71776 8236 71780
rect 8252 71836 8316 71840
rect 8252 71780 8256 71836
rect 8256 71780 8312 71836
rect 8312 71780 8316 71836
rect 8252 71776 8316 71780
rect 2352 71292 2416 71296
rect 2352 71236 2356 71292
rect 2356 71236 2412 71292
rect 2412 71236 2416 71292
rect 2352 71232 2416 71236
rect 2432 71292 2496 71296
rect 2432 71236 2436 71292
rect 2436 71236 2492 71292
rect 2492 71236 2496 71292
rect 2432 71232 2496 71236
rect 2512 71292 2576 71296
rect 2512 71236 2516 71292
rect 2516 71236 2572 71292
rect 2572 71236 2576 71292
rect 2512 71232 2576 71236
rect 2592 71292 2656 71296
rect 2592 71236 2596 71292
rect 2596 71236 2652 71292
rect 2652 71236 2656 71292
rect 2592 71232 2656 71236
rect 7352 71292 7416 71296
rect 7352 71236 7356 71292
rect 7356 71236 7412 71292
rect 7412 71236 7416 71292
rect 7352 71232 7416 71236
rect 7432 71292 7496 71296
rect 7432 71236 7436 71292
rect 7436 71236 7492 71292
rect 7492 71236 7496 71292
rect 7432 71232 7496 71236
rect 7512 71292 7576 71296
rect 7512 71236 7516 71292
rect 7516 71236 7572 71292
rect 7572 71236 7576 71292
rect 7512 71232 7576 71236
rect 7592 71292 7656 71296
rect 7592 71236 7596 71292
rect 7596 71236 7652 71292
rect 7652 71236 7656 71292
rect 7592 71232 7656 71236
rect 3012 70748 3076 70752
rect 3012 70692 3016 70748
rect 3016 70692 3072 70748
rect 3072 70692 3076 70748
rect 3012 70688 3076 70692
rect 3092 70748 3156 70752
rect 3092 70692 3096 70748
rect 3096 70692 3152 70748
rect 3152 70692 3156 70748
rect 3092 70688 3156 70692
rect 3172 70748 3236 70752
rect 3172 70692 3176 70748
rect 3176 70692 3232 70748
rect 3232 70692 3236 70748
rect 3172 70688 3236 70692
rect 3252 70748 3316 70752
rect 3252 70692 3256 70748
rect 3256 70692 3312 70748
rect 3312 70692 3316 70748
rect 3252 70688 3316 70692
rect 8012 70748 8076 70752
rect 8012 70692 8016 70748
rect 8016 70692 8072 70748
rect 8072 70692 8076 70748
rect 8012 70688 8076 70692
rect 8092 70748 8156 70752
rect 8092 70692 8096 70748
rect 8096 70692 8152 70748
rect 8152 70692 8156 70748
rect 8092 70688 8156 70692
rect 8172 70748 8236 70752
rect 8172 70692 8176 70748
rect 8176 70692 8232 70748
rect 8232 70692 8236 70748
rect 8172 70688 8236 70692
rect 8252 70748 8316 70752
rect 8252 70692 8256 70748
rect 8256 70692 8312 70748
rect 8312 70692 8316 70748
rect 8252 70688 8316 70692
rect 2352 70204 2416 70208
rect 2352 70148 2356 70204
rect 2356 70148 2412 70204
rect 2412 70148 2416 70204
rect 2352 70144 2416 70148
rect 2432 70204 2496 70208
rect 2432 70148 2436 70204
rect 2436 70148 2492 70204
rect 2492 70148 2496 70204
rect 2432 70144 2496 70148
rect 2512 70204 2576 70208
rect 2512 70148 2516 70204
rect 2516 70148 2572 70204
rect 2572 70148 2576 70204
rect 2512 70144 2576 70148
rect 2592 70204 2656 70208
rect 2592 70148 2596 70204
rect 2596 70148 2652 70204
rect 2652 70148 2656 70204
rect 2592 70144 2656 70148
rect 7352 70204 7416 70208
rect 7352 70148 7356 70204
rect 7356 70148 7412 70204
rect 7412 70148 7416 70204
rect 7352 70144 7416 70148
rect 7432 70204 7496 70208
rect 7432 70148 7436 70204
rect 7436 70148 7492 70204
rect 7492 70148 7496 70204
rect 7432 70144 7496 70148
rect 7512 70204 7576 70208
rect 7512 70148 7516 70204
rect 7516 70148 7572 70204
rect 7572 70148 7576 70204
rect 7512 70144 7576 70148
rect 7592 70204 7656 70208
rect 7592 70148 7596 70204
rect 7596 70148 7652 70204
rect 7652 70148 7656 70204
rect 7592 70144 7656 70148
rect 3012 69660 3076 69664
rect 3012 69604 3016 69660
rect 3016 69604 3072 69660
rect 3072 69604 3076 69660
rect 3012 69600 3076 69604
rect 3092 69660 3156 69664
rect 3092 69604 3096 69660
rect 3096 69604 3152 69660
rect 3152 69604 3156 69660
rect 3092 69600 3156 69604
rect 3172 69660 3236 69664
rect 3172 69604 3176 69660
rect 3176 69604 3232 69660
rect 3232 69604 3236 69660
rect 3172 69600 3236 69604
rect 3252 69660 3316 69664
rect 3252 69604 3256 69660
rect 3256 69604 3312 69660
rect 3312 69604 3316 69660
rect 3252 69600 3316 69604
rect 8012 69660 8076 69664
rect 8012 69604 8016 69660
rect 8016 69604 8072 69660
rect 8072 69604 8076 69660
rect 8012 69600 8076 69604
rect 8092 69660 8156 69664
rect 8092 69604 8096 69660
rect 8096 69604 8152 69660
rect 8152 69604 8156 69660
rect 8092 69600 8156 69604
rect 8172 69660 8236 69664
rect 8172 69604 8176 69660
rect 8176 69604 8232 69660
rect 8232 69604 8236 69660
rect 8172 69600 8236 69604
rect 8252 69660 8316 69664
rect 8252 69604 8256 69660
rect 8256 69604 8312 69660
rect 8312 69604 8316 69660
rect 8252 69600 8316 69604
rect 2352 69116 2416 69120
rect 2352 69060 2356 69116
rect 2356 69060 2412 69116
rect 2412 69060 2416 69116
rect 2352 69056 2416 69060
rect 2432 69116 2496 69120
rect 2432 69060 2436 69116
rect 2436 69060 2492 69116
rect 2492 69060 2496 69116
rect 2432 69056 2496 69060
rect 2512 69116 2576 69120
rect 2512 69060 2516 69116
rect 2516 69060 2572 69116
rect 2572 69060 2576 69116
rect 2512 69056 2576 69060
rect 2592 69116 2656 69120
rect 2592 69060 2596 69116
rect 2596 69060 2652 69116
rect 2652 69060 2656 69116
rect 2592 69056 2656 69060
rect 7352 69116 7416 69120
rect 7352 69060 7356 69116
rect 7356 69060 7412 69116
rect 7412 69060 7416 69116
rect 7352 69056 7416 69060
rect 7432 69116 7496 69120
rect 7432 69060 7436 69116
rect 7436 69060 7492 69116
rect 7492 69060 7496 69116
rect 7432 69056 7496 69060
rect 7512 69116 7576 69120
rect 7512 69060 7516 69116
rect 7516 69060 7572 69116
rect 7572 69060 7576 69116
rect 7512 69056 7576 69060
rect 7592 69116 7656 69120
rect 7592 69060 7596 69116
rect 7596 69060 7652 69116
rect 7652 69060 7656 69116
rect 7592 69056 7656 69060
rect 3012 68572 3076 68576
rect 3012 68516 3016 68572
rect 3016 68516 3072 68572
rect 3072 68516 3076 68572
rect 3012 68512 3076 68516
rect 3092 68572 3156 68576
rect 3092 68516 3096 68572
rect 3096 68516 3152 68572
rect 3152 68516 3156 68572
rect 3092 68512 3156 68516
rect 3172 68572 3236 68576
rect 3172 68516 3176 68572
rect 3176 68516 3232 68572
rect 3232 68516 3236 68572
rect 3172 68512 3236 68516
rect 3252 68572 3316 68576
rect 3252 68516 3256 68572
rect 3256 68516 3312 68572
rect 3312 68516 3316 68572
rect 3252 68512 3316 68516
rect 8012 68572 8076 68576
rect 8012 68516 8016 68572
rect 8016 68516 8072 68572
rect 8072 68516 8076 68572
rect 8012 68512 8076 68516
rect 8092 68572 8156 68576
rect 8092 68516 8096 68572
rect 8096 68516 8152 68572
rect 8152 68516 8156 68572
rect 8092 68512 8156 68516
rect 8172 68572 8236 68576
rect 8172 68516 8176 68572
rect 8176 68516 8232 68572
rect 8232 68516 8236 68572
rect 8172 68512 8236 68516
rect 8252 68572 8316 68576
rect 8252 68516 8256 68572
rect 8256 68516 8312 68572
rect 8312 68516 8316 68572
rect 8252 68512 8316 68516
rect 2352 68028 2416 68032
rect 2352 67972 2356 68028
rect 2356 67972 2412 68028
rect 2412 67972 2416 68028
rect 2352 67968 2416 67972
rect 2432 68028 2496 68032
rect 2432 67972 2436 68028
rect 2436 67972 2492 68028
rect 2492 67972 2496 68028
rect 2432 67968 2496 67972
rect 2512 68028 2576 68032
rect 2512 67972 2516 68028
rect 2516 67972 2572 68028
rect 2572 67972 2576 68028
rect 2512 67968 2576 67972
rect 2592 68028 2656 68032
rect 2592 67972 2596 68028
rect 2596 67972 2652 68028
rect 2652 67972 2656 68028
rect 2592 67968 2656 67972
rect 7352 68028 7416 68032
rect 7352 67972 7356 68028
rect 7356 67972 7412 68028
rect 7412 67972 7416 68028
rect 7352 67968 7416 67972
rect 7432 68028 7496 68032
rect 7432 67972 7436 68028
rect 7436 67972 7492 68028
rect 7492 67972 7496 68028
rect 7432 67968 7496 67972
rect 7512 68028 7576 68032
rect 7512 67972 7516 68028
rect 7516 67972 7572 68028
rect 7572 67972 7576 68028
rect 7512 67968 7576 67972
rect 7592 68028 7656 68032
rect 7592 67972 7596 68028
rect 7596 67972 7652 68028
rect 7652 67972 7656 68028
rect 7592 67968 7656 67972
rect 3012 67484 3076 67488
rect 3012 67428 3016 67484
rect 3016 67428 3072 67484
rect 3072 67428 3076 67484
rect 3012 67424 3076 67428
rect 3092 67484 3156 67488
rect 3092 67428 3096 67484
rect 3096 67428 3152 67484
rect 3152 67428 3156 67484
rect 3092 67424 3156 67428
rect 3172 67484 3236 67488
rect 3172 67428 3176 67484
rect 3176 67428 3232 67484
rect 3232 67428 3236 67484
rect 3172 67424 3236 67428
rect 3252 67484 3316 67488
rect 3252 67428 3256 67484
rect 3256 67428 3312 67484
rect 3312 67428 3316 67484
rect 3252 67424 3316 67428
rect 8012 67484 8076 67488
rect 8012 67428 8016 67484
rect 8016 67428 8072 67484
rect 8072 67428 8076 67484
rect 8012 67424 8076 67428
rect 8092 67484 8156 67488
rect 8092 67428 8096 67484
rect 8096 67428 8152 67484
rect 8152 67428 8156 67484
rect 8092 67424 8156 67428
rect 8172 67484 8236 67488
rect 8172 67428 8176 67484
rect 8176 67428 8232 67484
rect 8232 67428 8236 67484
rect 8172 67424 8236 67428
rect 8252 67484 8316 67488
rect 8252 67428 8256 67484
rect 8256 67428 8312 67484
rect 8312 67428 8316 67484
rect 8252 67424 8316 67428
rect 2352 66940 2416 66944
rect 2352 66884 2356 66940
rect 2356 66884 2412 66940
rect 2412 66884 2416 66940
rect 2352 66880 2416 66884
rect 2432 66940 2496 66944
rect 2432 66884 2436 66940
rect 2436 66884 2492 66940
rect 2492 66884 2496 66940
rect 2432 66880 2496 66884
rect 2512 66940 2576 66944
rect 2512 66884 2516 66940
rect 2516 66884 2572 66940
rect 2572 66884 2576 66940
rect 2512 66880 2576 66884
rect 2592 66940 2656 66944
rect 2592 66884 2596 66940
rect 2596 66884 2652 66940
rect 2652 66884 2656 66940
rect 2592 66880 2656 66884
rect 7352 66940 7416 66944
rect 7352 66884 7356 66940
rect 7356 66884 7412 66940
rect 7412 66884 7416 66940
rect 7352 66880 7416 66884
rect 7432 66940 7496 66944
rect 7432 66884 7436 66940
rect 7436 66884 7492 66940
rect 7492 66884 7496 66940
rect 7432 66880 7496 66884
rect 7512 66940 7576 66944
rect 7512 66884 7516 66940
rect 7516 66884 7572 66940
rect 7572 66884 7576 66940
rect 7512 66880 7576 66884
rect 7592 66940 7656 66944
rect 7592 66884 7596 66940
rect 7596 66884 7652 66940
rect 7652 66884 7656 66940
rect 7592 66880 7656 66884
rect 3012 66396 3076 66400
rect 3012 66340 3016 66396
rect 3016 66340 3072 66396
rect 3072 66340 3076 66396
rect 3012 66336 3076 66340
rect 3092 66396 3156 66400
rect 3092 66340 3096 66396
rect 3096 66340 3152 66396
rect 3152 66340 3156 66396
rect 3092 66336 3156 66340
rect 3172 66396 3236 66400
rect 3172 66340 3176 66396
rect 3176 66340 3232 66396
rect 3232 66340 3236 66396
rect 3172 66336 3236 66340
rect 3252 66396 3316 66400
rect 3252 66340 3256 66396
rect 3256 66340 3312 66396
rect 3312 66340 3316 66396
rect 3252 66336 3316 66340
rect 8012 66396 8076 66400
rect 8012 66340 8016 66396
rect 8016 66340 8072 66396
rect 8072 66340 8076 66396
rect 8012 66336 8076 66340
rect 8092 66396 8156 66400
rect 8092 66340 8096 66396
rect 8096 66340 8152 66396
rect 8152 66340 8156 66396
rect 8092 66336 8156 66340
rect 8172 66396 8236 66400
rect 8172 66340 8176 66396
rect 8176 66340 8232 66396
rect 8232 66340 8236 66396
rect 8172 66336 8236 66340
rect 8252 66396 8316 66400
rect 8252 66340 8256 66396
rect 8256 66340 8312 66396
rect 8312 66340 8316 66396
rect 8252 66336 8316 66340
rect 2352 65852 2416 65856
rect 2352 65796 2356 65852
rect 2356 65796 2412 65852
rect 2412 65796 2416 65852
rect 2352 65792 2416 65796
rect 2432 65852 2496 65856
rect 2432 65796 2436 65852
rect 2436 65796 2492 65852
rect 2492 65796 2496 65852
rect 2432 65792 2496 65796
rect 2512 65852 2576 65856
rect 2512 65796 2516 65852
rect 2516 65796 2572 65852
rect 2572 65796 2576 65852
rect 2512 65792 2576 65796
rect 2592 65852 2656 65856
rect 2592 65796 2596 65852
rect 2596 65796 2652 65852
rect 2652 65796 2656 65852
rect 2592 65792 2656 65796
rect 7352 65852 7416 65856
rect 7352 65796 7356 65852
rect 7356 65796 7412 65852
rect 7412 65796 7416 65852
rect 7352 65792 7416 65796
rect 7432 65852 7496 65856
rect 7432 65796 7436 65852
rect 7436 65796 7492 65852
rect 7492 65796 7496 65852
rect 7432 65792 7496 65796
rect 7512 65852 7576 65856
rect 7512 65796 7516 65852
rect 7516 65796 7572 65852
rect 7572 65796 7576 65852
rect 7512 65792 7576 65796
rect 7592 65852 7656 65856
rect 7592 65796 7596 65852
rect 7596 65796 7652 65852
rect 7652 65796 7656 65852
rect 7592 65792 7656 65796
rect 3012 65308 3076 65312
rect 3012 65252 3016 65308
rect 3016 65252 3072 65308
rect 3072 65252 3076 65308
rect 3012 65248 3076 65252
rect 3092 65308 3156 65312
rect 3092 65252 3096 65308
rect 3096 65252 3152 65308
rect 3152 65252 3156 65308
rect 3092 65248 3156 65252
rect 3172 65308 3236 65312
rect 3172 65252 3176 65308
rect 3176 65252 3232 65308
rect 3232 65252 3236 65308
rect 3172 65248 3236 65252
rect 3252 65308 3316 65312
rect 3252 65252 3256 65308
rect 3256 65252 3312 65308
rect 3312 65252 3316 65308
rect 3252 65248 3316 65252
rect 8012 65308 8076 65312
rect 8012 65252 8016 65308
rect 8016 65252 8072 65308
rect 8072 65252 8076 65308
rect 8012 65248 8076 65252
rect 8092 65308 8156 65312
rect 8092 65252 8096 65308
rect 8096 65252 8152 65308
rect 8152 65252 8156 65308
rect 8092 65248 8156 65252
rect 8172 65308 8236 65312
rect 8172 65252 8176 65308
rect 8176 65252 8232 65308
rect 8232 65252 8236 65308
rect 8172 65248 8236 65252
rect 8252 65308 8316 65312
rect 8252 65252 8256 65308
rect 8256 65252 8312 65308
rect 8312 65252 8316 65308
rect 8252 65248 8316 65252
rect 2352 64764 2416 64768
rect 2352 64708 2356 64764
rect 2356 64708 2412 64764
rect 2412 64708 2416 64764
rect 2352 64704 2416 64708
rect 2432 64764 2496 64768
rect 2432 64708 2436 64764
rect 2436 64708 2492 64764
rect 2492 64708 2496 64764
rect 2432 64704 2496 64708
rect 2512 64764 2576 64768
rect 2512 64708 2516 64764
rect 2516 64708 2572 64764
rect 2572 64708 2576 64764
rect 2512 64704 2576 64708
rect 2592 64764 2656 64768
rect 2592 64708 2596 64764
rect 2596 64708 2652 64764
rect 2652 64708 2656 64764
rect 2592 64704 2656 64708
rect 7352 64764 7416 64768
rect 7352 64708 7356 64764
rect 7356 64708 7412 64764
rect 7412 64708 7416 64764
rect 7352 64704 7416 64708
rect 7432 64764 7496 64768
rect 7432 64708 7436 64764
rect 7436 64708 7492 64764
rect 7492 64708 7496 64764
rect 7432 64704 7496 64708
rect 7512 64764 7576 64768
rect 7512 64708 7516 64764
rect 7516 64708 7572 64764
rect 7572 64708 7576 64764
rect 7512 64704 7576 64708
rect 7592 64764 7656 64768
rect 7592 64708 7596 64764
rect 7596 64708 7652 64764
rect 7652 64708 7656 64764
rect 7592 64704 7656 64708
rect 3012 64220 3076 64224
rect 3012 64164 3016 64220
rect 3016 64164 3072 64220
rect 3072 64164 3076 64220
rect 3012 64160 3076 64164
rect 3092 64220 3156 64224
rect 3092 64164 3096 64220
rect 3096 64164 3152 64220
rect 3152 64164 3156 64220
rect 3092 64160 3156 64164
rect 3172 64220 3236 64224
rect 3172 64164 3176 64220
rect 3176 64164 3232 64220
rect 3232 64164 3236 64220
rect 3172 64160 3236 64164
rect 3252 64220 3316 64224
rect 3252 64164 3256 64220
rect 3256 64164 3312 64220
rect 3312 64164 3316 64220
rect 3252 64160 3316 64164
rect 8012 64220 8076 64224
rect 8012 64164 8016 64220
rect 8016 64164 8072 64220
rect 8072 64164 8076 64220
rect 8012 64160 8076 64164
rect 8092 64220 8156 64224
rect 8092 64164 8096 64220
rect 8096 64164 8152 64220
rect 8152 64164 8156 64220
rect 8092 64160 8156 64164
rect 8172 64220 8236 64224
rect 8172 64164 8176 64220
rect 8176 64164 8232 64220
rect 8232 64164 8236 64220
rect 8172 64160 8236 64164
rect 8252 64220 8316 64224
rect 8252 64164 8256 64220
rect 8256 64164 8312 64220
rect 8312 64164 8316 64220
rect 8252 64160 8316 64164
rect 2352 63676 2416 63680
rect 2352 63620 2356 63676
rect 2356 63620 2412 63676
rect 2412 63620 2416 63676
rect 2352 63616 2416 63620
rect 2432 63676 2496 63680
rect 2432 63620 2436 63676
rect 2436 63620 2492 63676
rect 2492 63620 2496 63676
rect 2432 63616 2496 63620
rect 2512 63676 2576 63680
rect 2512 63620 2516 63676
rect 2516 63620 2572 63676
rect 2572 63620 2576 63676
rect 2512 63616 2576 63620
rect 2592 63676 2656 63680
rect 2592 63620 2596 63676
rect 2596 63620 2652 63676
rect 2652 63620 2656 63676
rect 2592 63616 2656 63620
rect 7352 63676 7416 63680
rect 7352 63620 7356 63676
rect 7356 63620 7412 63676
rect 7412 63620 7416 63676
rect 7352 63616 7416 63620
rect 7432 63676 7496 63680
rect 7432 63620 7436 63676
rect 7436 63620 7492 63676
rect 7492 63620 7496 63676
rect 7432 63616 7496 63620
rect 7512 63676 7576 63680
rect 7512 63620 7516 63676
rect 7516 63620 7572 63676
rect 7572 63620 7576 63676
rect 7512 63616 7576 63620
rect 7592 63676 7656 63680
rect 7592 63620 7596 63676
rect 7596 63620 7652 63676
rect 7652 63620 7656 63676
rect 7592 63616 7656 63620
rect 3012 63132 3076 63136
rect 3012 63076 3016 63132
rect 3016 63076 3072 63132
rect 3072 63076 3076 63132
rect 3012 63072 3076 63076
rect 3092 63132 3156 63136
rect 3092 63076 3096 63132
rect 3096 63076 3152 63132
rect 3152 63076 3156 63132
rect 3092 63072 3156 63076
rect 3172 63132 3236 63136
rect 3172 63076 3176 63132
rect 3176 63076 3232 63132
rect 3232 63076 3236 63132
rect 3172 63072 3236 63076
rect 3252 63132 3316 63136
rect 3252 63076 3256 63132
rect 3256 63076 3312 63132
rect 3312 63076 3316 63132
rect 3252 63072 3316 63076
rect 8012 63132 8076 63136
rect 8012 63076 8016 63132
rect 8016 63076 8072 63132
rect 8072 63076 8076 63132
rect 8012 63072 8076 63076
rect 8092 63132 8156 63136
rect 8092 63076 8096 63132
rect 8096 63076 8152 63132
rect 8152 63076 8156 63132
rect 8092 63072 8156 63076
rect 8172 63132 8236 63136
rect 8172 63076 8176 63132
rect 8176 63076 8232 63132
rect 8232 63076 8236 63132
rect 8172 63072 8236 63076
rect 8252 63132 8316 63136
rect 8252 63076 8256 63132
rect 8256 63076 8312 63132
rect 8312 63076 8316 63132
rect 8252 63072 8316 63076
rect 2352 62588 2416 62592
rect 2352 62532 2356 62588
rect 2356 62532 2412 62588
rect 2412 62532 2416 62588
rect 2352 62528 2416 62532
rect 2432 62588 2496 62592
rect 2432 62532 2436 62588
rect 2436 62532 2492 62588
rect 2492 62532 2496 62588
rect 2432 62528 2496 62532
rect 2512 62588 2576 62592
rect 2512 62532 2516 62588
rect 2516 62532 2572 62588
rect 2572 62532 2576 62588
rect 2512 62528 2576 62532
rect 2592 62588 2656 62592
rect 2592 62532 2596 62588
rect 2596 62532 2652 62588
rect 2652 62532 2656 62588
rect 2592 62528 2656 62532
rect 7352 62588 7416 62592
rect 7352 62532 7356 62588
rect 7356 62532 7412 62588
rect 7412 62532 7416 62588
rect 7352 62528 7416 62532
rect 7432 62588 7496 62592
rect 7432 62532 7436 62588
rect 7436 62532 7492 62588
rect 7492 62532 7496 62588
rect 7432 62528 7496 62532
rect 7512 62588 7576 62592
rect 7512 62532 7516 62588
rect 7516 62532 7572 62588
rect 7572 62532 7576 62588
rect 7512 62528 7576 62532
rect 7592 62588 7656 62592
rect 7592 62532 7596 62588
rect 7596 62532 7652 62588
rect 7652 62532 7656 62588
rect 7592 62528 7656 62532
rect 3012 62044 3076 62048
rect 3012 61988 3016 62044
rect 3016 61988 3072 62044
rect 3072 61988 3076 62044
rect 3012 61984 3076 61988
rect 3092 62044 3156 62048
rect 3092 61988 3096 62044
rect 3096 61988 3152 62044
rect 3152 61988 3156 62044
rect 3092 61984 3156 61988
rect 3172 62044 3236 62048
rect 3172 61988 3176 62044
rect 3176 61988 3232 62044
rect 3232 61988 3236 62044
rect 3172 61984 3236 61988
rect 3252 62044 3316 62048
rect 3252 61988 3256 62044
rect 3256 61988 3312 62044
rect 3312 61988 3316 62044
rect 3252 61984 3316 61988
rect 8012 62044 8076 62048
rect 8012 61988 8016 62044
rect 8016 61988 8072 62044
rect 8072 61988 8076 62044
rect 8012 61984 8076 61988
rect 8092 62044 8156 62048
rect 8092 61988 8096 62044
rect 8096 61988 8152 62044
rect 8152 61988 8156 62044
rect 8092 61984 8156 61988
rect 8172 62044 8236 62048
rect 8172 61988 8176 62044
rect 8176 61988 8232 62044
rect 8232 61988 8236 62044
rect 8172 61984 8236 61988
rect 8252 62044 8316 62048
rect 8252 61988 8256 62044
rect 8256 61988 8312 62044
rect 8312 61988 8316 62044
rect 8252 61984 8316 61988
rect 2352 61500 2416 61504
rect 2352 61444 2356 61500
rect 2356 61444 2412 61500
rect 2412 61444 2416 61500
rect 2352 61440 2416 61444
rect 2432 61500 2496 61504
rect 2432 61444 2436 61500
rect 2436 61444 2492 61500
rect 2492 61444 2496 61500
rect 2432 61440 2496 61444
rect 2512 61500 2576 61504
rect 2512 61444 2516 61500
rect 2516 61444 2572 61500
rect 2572 61444 2576 61500
rect 2512 61440 2576 61444
rect 2592 61500 2656 61504
rect 2592 61444 2596 61500
rect 2596 61444 2652 61500
rect 2652 61444 2656 61500
rect 2592 61440 2656 61444
rect 7352 61500 7416 61504
rect 7352 61444 7356 61500
rect 7356 61444 7412 61500
rect 7412 61444 7416 61500
rect 7352 61440 7416 61444
rect 7432 61500 7496 61504
rect 7432 61444 7436 61500
rect 7436 61444 7492 61500
rect 7492 61444 7496 61500
rect 7432 61440 7496 61444
rect 7512 61500 7576 61504
rect 7512 61444 7516 61500
rect 7516 61444 7572 61500
rect 7572 61444 7576 61500
rect 7512 61440 7576 61444
rect 7592 61500 7656 61504
rect 7592 61444 7596 61500
rect 7596 61444 7652 61500
rect 7652 61444 7656 61500
rect 7592 61440 7656 61444
rect 3012 60956 3076 60960
rect 3012 60900 3016 60956
rect 3016 60900 3072 60956
rect 3072 60900 3076 60956
rect 3012 60896 3076 60900
rect 3092 60956 3156 60960
rect 3092 60900 3096 60956
rect 3096 60900 3152 60956
rect 3152 60900 3156 60956
rect 3092 60896 3156 60900
rect 3172 60956 3236 60960
rect 3172 60900 3176 60956
rect 3176 60900 3232 60956
rect 3232 60900 3236 60956
rect 3172 60896 3236 60900
rect 3252 60956 3316 60960
rect 3252 60900 3256 60956
rect 3256 60900 3312 60956
rect 3312 60900 3316 60956
rect 3252 60896 3316 60900
rect 8012 60956 8076 60960
rect 8012 60900 8016 60956
rect 8016 60900 8072 60956
rect 8072 60900 8076 60956
rect 8012 60896 8076 60900
rect 8092 60956 8156 60960
rect 8092 60900 8096 60956
rect 8096 60900 8152 60956
rect 8152 60900 8156 60956
rect 8092 60896 8156 60900
rect 8172 60956 8236 60960
rect 8172 60900 8176 60956
rect 8176 60900 8232 60956
rect 8232 60900 8236 60956
rect 8172 60896 8236 60900
rect 8252 60956 8316 60960
rect 8252 60900 8256 60956
rect 8256 60900 8312 60956
rect 8312 60900 8316 60956
rect 8252 60896 8316 60900
rect 2352 60412 2416 60416
rect 2352 60356 2356 60412
rect 2356 60356 2412 60412
rect 2412 60356 2416 60412
rect 2352 60352 2416 60356
rect 2432 60412 2496 60416
rect 2432 60356 2436 60412
rect 2436 60356 2492 60412
rect 2492 60356 2496 60412
rect 2432 60352 2496 60356
rect 2512 60412 2576 60416
rect 2512 60356 2516 60412
rect 2516 60356 2572 60412
rect 2572 60356 2576 60412
rect 2512 60352 2576 60356
rect 2592 60412 2656 60416
rect 2592 60356 2596 60412
rect 2596 60356 2652 60412
rect 2652 60356 2656 60412
rect 2592 60352 2656 60356
rect 7352 60412 7416 60416
rect 7352 60356 7356 60412
rect 7356 60356 7412 60412
rect 7412 60356 7416 60412
rect 7352 60352 7416 60356
rect 7432 60412 7496 60416
rect 7432 60356 7436 60412
rect 7436 60356 7492 60412
rect 7492 60356 7496 60412
rect 7432 60352 7496 60356
rect 7512 60412 7576 60416
rect 7512 60356 7516 60412
rect 7516 60356 7572 60412
rect 7572 60356 7576 60412
rect 7512 60352 7576 60356
rect 7592 60412 7656 60416
rect 7592 60356 7596 60412
rect 7596 60356 7652 60412
rect 7652 60356 7656 60412
rect 7592 60352 7656 60356
rect 3012 59868 3076 59872
rect 3012 59812 3016 59868
rect 3016 59812 3072 59868
rect 3072 59812 3076 59868
rect 3012 59808 3076 59812
rect 3092 59868 3156 59872
rect 3092 59812 3096 59868
rect 3096 59812 3152 59868
rect 3152 59812 3156 59868
rect 3092 59808 3156 59812
rect 3172 59868 3236 59872
rect 3172 59812 3176 59868
rect 3176 59812 3232 59868
rect 3232 59812 3236 59868
rect 3172 59808 3236 59812
rect 3252 59868 3316 59872
rect 3252 59812 3256 59868
rect 3256 59812 3312 59868
rect 3312 59812 3316 59868
rect 3252 59808 3316 59812
rect 8012 59868 8076 59872
rect 8012 59812 8016 59868
rect 8016 59812 8072 59868
rect 8072 59812 8076 59868
rect 8012 59808 8076 59812
rect 8092 59868 8156 59872
rect 8092 59812 8096 59868
rect 8096 59812 8152 59868
rect 8152 59812 8156 59868
rect 8092 59808 8156 59812
rect 8172 59868 8236 59872
rect 8172 59812 8176 59868
rect 8176 59812 8232 59868
rect 8232 59812 8236 59868
rect 8172 59808 8236 59812
rect 8252 59868 8316 59872
rect 8252 59812 8256 59868
rect 8256 59812 8312 59868
rect 8312 59812 8316 59868
rect 8252 59808 8316 59812
rect 2352 59324 2416 59328
rect 2352 59268 2356 59324
rect 2356 59268 2412 59324
rect 2412 59268 2416 59324
rect 2352 59264 2416 59268
rect 2432 59324 2496 59328
rect 2432 59268 2436 59324
rect 2436 59268 2492 59324
rect 2492 59268 2496 59324
rect 2432 59264 2496 59268
rect 2512 59324 2576 59328
rect 2512 59268 2516 59324
rect 2516 59268 2572 59324
rect 2572 59268 2576 59324
rect 2512 59264 2576 59268
rect 2592 59324 2656 59328
rect 2592 59268 2596 59324
rect 2596 59268 2652 59324
rect 2652 59268 2656 59324
rect 2592 59264 2656 59268
rect 7352 59324 7416 59328
rect 7352 59268 7356 59324
rect 7356 59268 7412 59324
rect 7412 59268 7416 59324
rect 7352 59264 7416 59268
rect 7432 59324 7496 59328
rect 7432 59268 7436 59324
rect 7436 59268 7492 59324
rect 7492 59268 7496 59324
rect 7432 59264 7496 59268
rect 7512 59324 7576 59328
rect 7512 59268 7516 59324
rect 7516 59268 7572 59324
rect 7572 59268 7576 59324
rect 7512 59264 7576 59268
rect 7592 59324 7656 59328
rect 7592 59268 7596 59324
rect 7596 59268 7652 59324
rect 7652 59268 7656 59324
rect 7592 59264 7656 59268
rect 3012 58780 3076 58784
rect 3012 58724 3016 58780
rect 3016 58724 3072 58780
rect 3072 58724 3076 58780
rect 3012 58720 3076 58724
rect 3092 58780 3156 58784
rect 3092 58724 3096 58780
rect 3096 58724 3152 58780
rect 3152 58724 3156 58780
rect 3092 58720 3156 58724
rect 3172 58780 3236 58784
rect 3172 58724 3176 58780
rect 3176 58724 3232 58780
rect 3232 58724 3236 58780
rect 3172 58720 3236 58724
rect 3252 58780 3316 58784
rect 3252 58724 3256 58780
rect 3256 58724 3312 58780
rect 3312 58724 3316 58780
rect 3252 58720 3316 58724
rect 8012 58780 8076 58784
rect 8012 58724 8016 58780
rect 8016 58724 8072 58780
rect 8072 58724 8076 58780
rect 8012 58720 8076 58724
rect 8092 58780 8156 58784
rect 8092 58724 8096 58780
rect 8096 58724 8152 58780
rect 8152 58724 8156 58780
rect 8092 58720 8156 58724
rect 8172 58780 8236 58784
rect 8172 58724 8176 58780
rect 8176 58724 8232 58780
rect 8232 58724 8236 58780
rect 8172 58720 8236 58724
rect 8252 58780 8316 58784
rect 8252 58724 8256 58780
rect 8256 58724 8312 58780
rect 8312 58724 8316 58780
rect 8252 58720 8316 58724
rect 2352 58236 2416 58240
rect 2352 58180 2356 58236
rect 2356 58180 2412 58236
rect 2412 58180 2416 58236
rect 2352 58176 2416 58180
rect 2432 58236 2496 58240
rect 2432 58180 2436 58236
rect 2436 58180 2492 58236
rect 2492 58180 2496 58236
rect 2432 58176 2496 58180
rect 2512 58236 2576 58240
rect 2512 58180 2516 58236
rect 2516 58180 2572 58236
rect 2572 58180 2576 58236
rect 2512 58176 2576 58180
rect 2592 58236 2656 58240
rect 2592 58180 2596 58236
rect 2596 58180 2652 58236
rect 2652 58180 2656 58236
rect 2592 58176 2656 58180
rect 7352 58236 7416 58240
rect 7352 58180 7356 58236
rect 7356 58180 7412 58236
rect 7412 58180 7416 58236
rect 7352 58176 7416 58180
rect 7432 58236 7496 58240
rect 7432 58180 7436 58236
rect 7436 58180 7492 58236
rect 7492 58180 7496 58236
rect 7432 58176 7496 58180
rect 7512 58236 7576 58240
rect 7512 58180 7516 58236
rect 7516 58180 7572 58236
rect 7572 58180 7576 58236
rect 7512 58176 7576 58180
rect 7592 58236 7656 58240
rect 7592 58180 7596 58236
rect 7596 58180 7652 58236
rect 7652 58180 7656 58236
rect 7592 58176 7656 58180
rect 3012 57692 3076 57696
rect 3012 57636 3016 57692
rect 3016 57636 3072 57692
rect 3072 57636 3076 57692
rect 3012 57632 3076 57636
rect 3092 57692 3156 57696
rect 3092 57636 3096 57692
rect 3096 57636 3152 57692
rect 3152 57636 3156 57692
rect 3092 57632 3156 57636
rect 3172 57692 3236 57696
rect 3172 57636 3176 57692
rect 3176 57636 3232 57692
rect 3232 57636 3236 57692
rect 3172 57632 3236 57636
rect 3252 57692 3316 57696
rect 3252 57636 3256 57692
rect 3256 57636 3312 57692
rect 3312 57636 3316 57692
rect 3252 57632 3316 57636
rect 8012 57692 8076 57696
rect 8012 57636 8016 57692
rect 8016 57636 8072 57692
rect 8072 57636 8076 57692
rect 8012 57632 8076 57636
rect 8092 57692 8156 57696
rect 8092 57636 8096 57692
rect 8096 57636 8152 57692
rect 8152 57636 8156 57692
rect 8092 57632 8156 57636
rect 8172 57692 8236 57696
rect 8172 57636 8176 57692
rect 8176 57636 8232 57692
rect 8232 57636 8236 57692
rect 8172 57632 8236 57636
rect 8252 57692 8316 57696
rect 8252 57636 8256 57692
rect 8256 57636 8312 57692
rect 8312 57636 8316 57692
rect 8252 57632 8316 57636
rect 2352 57148 2416 57152
rect 2352 57092 2356 57148
rect 2356 57092 2412 57148
rect 2412 57092 2416 57148
rect 2352 57088 2416 57092
rect 2432 57148 2496 57152
rect 2432 57092 2436 57148
rect 2436 57092 2492 57148
rect 2492 57092 2496 57148
rect 2432 57088 2496 57092
rect 2512 57148 2576 57152
rect 2512 57092 2516 57148
rect 2516 57092 2572 57148
rect 2572 57092 2576 57148
rect 2512 57088 2576 57092
rect 2592 57148 2656 57152
rect 2592 57092 2596 57148
rect 2596 57092 2652 57148
rect 2652 57092 2656 57148
rect 2592 57088 2656 57092
rect 7352 57148 7416 57152
rect 7352 57092 7356 57148
rect 7356 57092 7412 57148
rect 7412 57092 7416 57148
rect 7352 57088 7416 57092
rect 7432 57148 7496 57152
rect 7432 57092 7436 57148
rect 7436 57092 7492 57148
rect 7492 57092 7496 57148
rect 7432 57088 7496 57092
rect 7512 57148 7576 57152
rect 7512 57092 7516 57148
rect 7516 57092 7572 57148
rect 7572 57092 7576 57148
rect 7512 57088 7576 57092
rect 7592 57148 7656 57152
rect 7592 57092 7596 57148
rect 7596 57092 7652 57148
rect 7652 57092 7656 57148
rect 7592 57088 7656 57092
rect 3012 56604 3076 56608
rect 3012 56548 3016 56604
rect 3016 56548 3072 56604
rect 3072 56548 3076 56604
rect 3012 56544 3076 56548
rect 3092 56604 3156 56608
rect 3092 56548 3096 56604
rect 3096 56548 3152 56604
rect 3152 56548 3156 56604
rect 3092 56544 3156 56548
rect 3172 56604 3236 56608
rect 3172 56548 3176 56604
rect 3176 56548 3232 56604
rect 3232 56548 3236 56604
rect 3172 56544 3236 56548
rect 3252 56604 3316 56608
rect 3252 56548 3256 56604
rect 3256 56548 3312 56604
rect 3312 56548 3316 56604
rect 3252 56544 3316 56548
rect 8012 56604 8076 56608
rect 8012 56548 8016 56604
rect 8016 56548 8072 56604
rect 8072 56548 8076 56604
rect 8012 56544 8076 56548
rect 8092 56604 8156 56608
rect 8092 56548 8096 56604
rect 8096 56548 8152 56604
rect 8152 56548 8156 56604
rect 8092 56544 8156 56548
rect 8172 56604 8236 56608
rect 8172 56548 8176 56604
rect 8176 56548 8232 56604
rect 8232 56548 8236 56604
rect 8172 56544 8236 56548
rect 8252 56604 8316 56608
rect 8252 56548 8256 56604
rect 8256 56548 8312 56604
rect 8312 56548 8316 56604
rect 8252 56544 8316 56548
rect 2352 56060 2416 56064
rect 2352 56004 2356 56060
rect 2356 56004 2412 56060
rect 2412 56004 2416 56060
rect 2352 56000 2416 56004
rect 2432 56060 2496 56064
rect 2432 56004 2436 56060
rect 2436 56004 2492 56060
rect 2492 56004 2496 56060
rect 2432 56000 2496 56004
rect 2512 56060 2576 56064
rect 2512 56004 2516 56060
rect 2516 56004 2572 56060
rect 2572 56004 2576 56060
rect 2512 56000 2576 56004
rect 2592 56060 2656 56064
rect 2592 56004 2596 56060
rect 2596 56004 2652 56060
rect 2652 56004 2656 56060
rect 2592 56000 2656 56004
rect 7352 56060 7416 56064
rect 7352 56004 7356 56060
rect 7356 56004 7412 56060
rect 7412 56004 7416 56060
rect 7352 56000 7416 56004
rect 7432 56060 7496 56064
rect 7432 56004 7436 56060
rect 7436 56004 7492 56060
rect 7492 56004 7496 56060
rect 7432 56000 7496 56004
rect 7512 56060 7576 56064
rect 7512 56004 7516 56060
rect 7516 56004 7572 56060
rect 7572 56004 7576 56060
rect 7512 56000 7576 56004
rect 7592 56060 7656 56064
rect 7592 56004 7596 56060
rect 7596 56004 7652 56060
rect 7652 56004 7656 56060
rect 7592 56000 7656 56004
rect 3012 55516 3076 55520
rect 3012 55460 3016 55516
rect 3016 55460 3072 55516
rect 3072 55460 3076 55516
rect 3012 55456 3076 55460
rect 3092 55516 3156 55520
rect 3092 55460 3096 55516
rect 3096 55460 3152 55516
rect 3152 55460 3156 55516
rect 3092 55456 3156 55460
rect 3172 55516 3236 55520
rect 3172 55460 3176 55516
rect 3176 55460 3232 55516
rect 3232 55460 3236 55516
rect 3172 55456 3236 55460
rect 3252 55516 3316 55520
rect 3252 55460 3256 55516
rect 3256 55460 3312 55516
rect 3312 55460 3316 55516
rect 3252 55456 3316 55460
rect 8012 55516 8076 55520
rect 8012 55460 8016 55516
rect 8016 55460 8072 55516
rect 8072 55460 8076 55516
rect 8012 55456 8076 55460
rect 8092 55516 8156 55520
rect 8092 55460 8096 55516
rect 8096 55460 8152 55516
rect 8152 55460 8156 55516
rect 8092 55456 8156 55460
rect 8172 55516 8236 55520
rect 8172 55460 8176 55516
rect 8176 55460 8232 55516
rect 8232 55460 8236 55516
rect 8172 55456 8236 55460
rect 8252 55516 8316 55520
rect 8252 55460 8256 55516
rect 8256 55460 8312 55516
rect 8312 55460 8316 55516
rect 8252 55456 8316 55460
rect 2352 54972 2416 54976
rect 2352 54916 2356 54972
rect 2356 54916 2412 54972
rect 2412 54916 2416 54972
rect 2352 54912 2416 54916
rect 2432 54972 2496 54976
rect 2432 54916 2436 54972
rect 2436 54916 2492 54972
rect 2492 54916 2496 54972
rect 2432 54912 2496 54916
rect 2512 54972 2576 54976
rect 2512 54916 2516 54972
rect 2516 54916 2572 54972
rect 2572 54916 2576 54972
rect 2512 54912 2576 54916
rect 2592 54972 2656 54976
rect 2592 54916 2596 54972
rect 2596 54916 2652 54972
rect 2652 54916 2656 54972
rect 2592 54912 2656 54916
rect 7352 54972 7416 54976
rect 7352 54916 7356 54972
rect 7356 54916 7412 54972
rect 7412 54916 7416 54972
rect 7352 54912 7416 54916
rect 7432 54972 7496 54976
rect 7432 54916 7436 54972
rect 7436 54916 7492 54972
rect 7492 54916 7496 54972
rect 7432 54912 7496 54916
rect 7512 54972 7576 54976
rect 7512 54916 7516 54972
rect 7516 54916 7572 54972
rect 7572 54916 7576 54972
rect 7512 54912 7576 54916
rect 7592 54972 7656 54976
rect 7592 54916 7596 54972
rect 7596 54916 7652 54972
rect 7652 54916 7656 54972
rect 7592 54912 7656 54916
rect 3012 54428 3076 54432
rect 3012 54372 3016 54428
rect 3016 54372 3072 54428
rect 3072 54372 3076 54428
rect 3012 54368 3076 54372
rect 3092 54428 3156 54432
rect 3092 54372 3096 54428
rect 3096 54372 3152 54428
rect 3152 54372 3156 54428
rect 3092 54368 3156 54372
rect 3172 54428 3236 54432
rect 3172 54372 3176 54428
rect 3176 54372 3232 54428
rect 3232 54372 3236 54428
rect 3172 54368 3236 54372
rect 3252 54428 3316 54432
rect 3252 54372 3256 54428
rect 3256 54372 3312 54428
rect 3312 54372 3316 54428
rect 3252 54368 3316 54372
rect 8012 54428 8076 54432
rect 8012 54372 8016 54428
rect 8016 54372 8072 54428
rect 8072 54372 8076 54428
rect 8012 54368 8076 54372
rect 8092 54428 8156 54432
rect 8092 54372 8096 54428
rect 8096 54372 8152 54428
rect 8152 54372 8156 54428
rect 8092 54368 8156 54372
rect 8172 54428 8236 54432
rect 8172 54372 8176 54428
rect 8176 54372 8232 54428
rect 8232 54372 8236 54428
rect 8172 54368 8236 54372
rect 8252 54428 8316 54432
rect 8252 54372 8256 54428
rect 8256 54372 8312 54428
rect 8312 54372 8316 54428
rect 8252 54368 8316 54372
rect 2352 53884 2416 53888
rect 2352 53828 2356 53884
rect 2356 53828 2412 53884
rect 2412 53828 2416 53884
rect 2352 53824 2416 53828
rect 2432 53884 2496 53888
rect 2432 53828 2436 53884
rect 2436 53828 2492 53884
rect 2492 53828 2496 53884
rect 2432 53824 2496 53828
rect 2512 53884 2576 53888
rect 2512 53828 2516 53884
rect 2516 53828 2572 53884
rect 2572 53828 2576 53884
rect 2512 53824 2576 53828
rect 2592 53884 2656 53888
rect 2592 53828 2596 53884
rect 2596 53828 2652 53884
rect 2652 53828 2656 53884
rect 2592 53824 2656 53828
rect 7352 53884 7416 53888
rect 7352 53828 7356 53884
rect 7356 53828 7412 53884
rect 7412 53828 7416 53884
rect 7352 53824 7416 53828
rect 7432 53884 7496 53888
rect 7432 53828 7436 53884
rect 7436 53828 7492 53884
rect 7492 53828 7496 53884
rect 7432 53824 7496 53828
rect 7512 53884 7576 53888
rect 7512 53828 7516 53884
rect 7516 53828 7572 53884
rect 7572 53828 7576 53884
rect 7512 53824 7576 53828
rect 7592 53884 7656 53888
rect 7592 53828 7596 53884
rect 7596 53828 7652 53884
rect 7652 53828 7656 53884
rect 7592 53824 7656 53828
rect 3012 53340 3076 53344
rect 3012 53284 3016 53340
rect 3016 53284 3072 53340
rect 3072 53284 3076 53340
rect 3012 53280 3076 53284
rect 3092 53340 3156 53344
rect 3092 53284 3096 53340
rect 3096 53284 3152 53340
rect 3152 53284 3156 53340
rect 3092 53280 3156 53284
rect 3172 53340 3236 53344
rect 3172 53284 3176 53340
rect 3176 53284 3232 53340
rect 3232 53284 3236 53340
rect 3172 53280 3236 53284
rect 3252 53340 3316 53344
rect 3252 53284 3256 53340
rect 3256 53284 3312 53340
rect 3312 53284 3316 53340
rect 3252 53280 3316 53284
rect 8012 53340 8076 53344
rect 8012 53284 8016 53340
rect 8016 53284 8072 53340
rect 8072 53284 8076 53340
rect 8012 53280 8076 53284
rect 8092 53340 8156 53344
rect 8092 53284 8096 53340
rect 8096 53284 8152 53340
rect 8152 53284 8156 53340
rect 8092 53280 8156 53284
rect 8172 53340 8236 53344
rect 8172 53284 8176 53340
rect 8176 53284 8232 53340
rect 8232 53284 8236 53340
rect 8172 53280 8236 53284
rect 8252 53340 8316 53344
rect 8252 53284 8256 53340
rect 8256 53284 8312 53340
rect 8312 53284 8316 53340
rect 8252 53280 8316 53284
rect 2352 52796 2416 52800
rect 2352 52740 2356 52796
rect 2356 52740 2412 52796
rect 2412 52740 2416 52796
rect 2352 52736 2416 52740
rect 2432 52796 2496 52800
rect 2432 52740 2436 52796
rect 2436 52740 2492 52796
rect 2492 52740 2496 52796
rect 2432 52736 2496 52740
rect 2512 52796 2576 52800
rect 2512 52740 2516 52796
rect 2516 52740 2572 52796
rect 2572 52740 2576 52796
rect 2512 52736 2576 52740
rect 2592 52796 2656 52800
rect 2592 52740 2596 52796
rect 2596 52740 2652 52796
rect 2652 52740 2656 52796
rect 2592 52736 2656 52740
rect 7352 52796 7416 52800
rect 7352 52740 7356 52796
rect 7356 52740 7412 52796
rect 7412 52740 7416 52796
rect 7352 52736 7416 52740
rect 7432 52796 7496 52800
rect 7432 52740 7436 52796
rect 7436 52740 7492 52796
rect 7492 52740 7496 52796
rect 7432 52736 7496 52740
rect 7512 52796 7576 52800
rect 7512 52740 7516 52796
rect 7516 52740 7572 52796
rect 7572 52740 7576 52796
rect 7512 52736 7576 52740
rect 7592 52796 7656 52800
rect 7592 52740 7596 52796
rect 7596 52740 7652 52796
rect 7652 52740 7656 52796
rect 7592 52736 7656 52740
rect 3012 52252 3076 52256
rect 3012 52196 3016 52252
rect 3016 52196 3072 52252
rect 3072 52196 3076 52252
rect 3012 52192 3076 52196
rect 3092 52252 3156 52256
rect 3092 52196 3096 52252
rect 3096 52196 3152 52252
rect 3152 52196 3156 52252
rect 3092 52192 3156 52196
rect 3172 52252 3236 52256
rect 3172 52196 3176 52252
rect 3176 52196 3232 52252
rect 3232 52196 3236 52252
rect 3172 52192 3236 52196
rect 3252 52252 3316 52256
rect 3252 52196 3256 52252
rect 3256 52196 3312 52252
rect 3312 52196 3316 52252
rect 3252 52192 3316 52196
rect 8012 52252 8076 52256
rect 8012 52196 8016 52252
rect 8016 52196 8072 52252
rect 8072 52196 8076 52252
rect 8012 52192 8076 52196
rect 8092 52252 8156 52256
rect 8092 52196 8096 52252
rect 8096 52196 8152 52252
rect 8152 52196 8156 52252
rect 8092 52192 8156 52196
rect 8172 52252 8236 52256
rect 8172 52196 8176 52252
rect 8176 52196 8232 52252
rect 8232 52196 8236 52252
rect 8172 52192 8236 52196
rect 8252 52252 8316 52256
rect 8252 52196 8256 52252
rect 8256 52196 8312 52252
rect 8312 52196 8316 52252
rect 8252 52192 8316 52196
rect 2352 51708 2416 51712
rect 2352 51652 2356 51708
rect 2356 51652 2412 51708
rect 2412 51652 2416 51708
rect 2352 51648 2416 51652
rect 2432 51708 2496 51712
rect 2432 51652 2436 51708
rect 2436 51652 2492 51708
rect 2492 51652 2496 51708
rect 2432 51648 2496 51652
rect 2512 51708 2576 51712
rect 2512 51652 2516 51708
rect 2516 51652 2572 51708
rect 2572 51652 2576 51708
rect 2512 51648 2576 51652
rect 2592 51708 2656 51712
rect 2592 51652 2596 51708
rect 2596 51652 2652 51708
rect 2652 51652 2656 51708
rect 2592 51648 2656 51652
rect 7352 51708 7416 51712
rect 7352 51652 7356 51708
rect 7356 51652 7412 51708
rect 7412 51652 7416 51708
rect 7352 51648 7416 51652
rect 7432 51708 7496 51712
rect 7432 51652 7436 51708
rect 7436 51652 7492 51708
rect 7492 51652 7496 51708
rect 7432 51648 7496 51652
rect 7512 51708 7576 51712
rect 7512 51652 7516 51708
rect 7516 51652 7572 51708
rect 7572 51652 7576 51708
rect 7512 51648 7576 51652
rect 7592 51708 7656 51712
rect 7592 51652 7596 51708
rect 7596 51652 7652 51708
rect 7652 51652 7656 51708
rect 7592 51648 7656 51652
rect 3012 51164 3076 51168
rect 3012 51108 3016 51164
rect 3016 51108 3072 51164
rect 3072 51108 3076 51164
rect 3012 51104 3076 51108
rect 3092 51164 3156 51168
rect 3092 51108 3096 51164
rect 3096 51108 3152 51164
rect 3152 51108 3156 51164
rect 3092 51104 3156 51108
rect 3172 51164 3236 51168
rect 3172 51108 3176 51164
rect 3176 51108 3232 51164
rect 3232 51108 3236 51164
rect 3172 51104 3236 51108
rect 3252 51164 3316 51168
rect 3252 51108 3256 51164
rect 3256 51108 3312 51164
rect 3312 51108 3316 51164
rect 3252 51104 3316 51108
rect 8012 51164 8076 51168
rect 8012 51108 8016 51164
rect 8016 51108 8072 51164
rect 8072 51108 8076 51164
rect 8012 51104 8076 51108
rect 8092 51164 8156 51168
rect 8092 51108 8096 51164
rect 8096 51108 8152 51164
rect 8152 51108 8156 51164
rect 8092 51104 8156 51108
rect 8172 51164 8236 51168
rect 8172 51108 8176 51164
rect 8176 51108 8232 51164
rect 8232 51108 8236 51164
rect 8172 51104 8236 51108
rect 8252 51164 8316 51168
rect 8252 51108 8256 51164
rect 8256 51108 8312 51164
rect 8312 51108 8316 51164
rect 8252 51104 8316 51108
rect 2352 50620 2416 50624
rect 2352 50564 2356 50620
rect 2356 50564 2412 50620
rect 2412 50564 2416 50620
rect 2352 50560 2416 50564
rect 2432 50620 2496 50624
rect 2432 50564 2436 50620
rect 2436 50564 2492 50620
rect 2492 50564 2496 50620
rect 2432 50560 2496 50564
rect 2512 50620 2576 50624
rect 2512 50564 2516 50620
rect 2516 50564 2572 50620
rect 2572 50564 2576 50620
rect 2512 50560 2576 50564
rect 2592 50620 2656 50624
rect 2592 50564 2596 50620
rect 2596 50564 2652 50620
rect 2652 50564 2656 50620
rect 2592 50560 2656 50564
rect 7352 50620 7416 50624
rect 7352 50564 7356 50620
rect 7356 50564 7412 50620
rect 7412 50564 7416 50620
rect 7352 50560 7416 50564
rect 7432 50620 7496 50624
rect 7432 50564 7436 50620
rect 7436 50564 7492 50620
rect 7492 50564 7496 50620
rect 7432 50560 7496 50564
rect 7512 50620 7576 50624
rect 7512 50564 7516 50620
rect 7516 50564 7572 50620
rect 7572 50564 7576 50620
rect 7512 50560 7576 50564
rect 7592 50620 7656 50624
rect 7592 50564 7596 50620
rect 7596 50564 7652 50620
rect 7652 50564 7656 50620
rect 7592 50560 7656 50564
rect 3012 50076 3076 50080
rect 3012 50020 3016 50076
rect 3016 50020 3072 50076
rect 3072 50020 3076 50076
rect 3012 50016 3076 50020
rect 3092 50076 3156 50080
rect 3092 50020 3096 50076
rect 3096 50020 3152 50076
rect 3152 50020 3156 50076
rect 3092 50016 3156 50020
rect 3172 50076 3236 50080
rect 3172 50020 3176 50076
rect 3176 50020 3232 50076
rect 3232 50020 3236 50076
rect 3172 50016 3236 50020
rect 3252 50076 3316 50080
rect 3252 50020 3256 50076
rect 3256 50020 3312 50076
rect 3312 50020 3316 50076
rect 3252 50016 3316 50020
rect 8012 50076 8076 50080
rect 8012 50020 8016 50076
rect 8016 50020 8072 50076
rect 8072 50020 8076 50076
rect 8012 50016 8076 50020
rect 8092 50076 8156 50080
rect 8092 50020 8096 50076
rect 8096 50020 8152 50076
rect 8152 50020 8156 50076
rect 8092 50016 8156 50020
rect 8172 50076 8236 50080
rect 8172 50020 8176 50076
rect 8176 50020 8232 50076
rect 8232 50020 8236 50076
rect 8172 50016 8236 50020
rect 8252 50076 8316 50080
rect 8252 50020 8256 50076
rect 8256 50020 8312 50076
rect 8312 50020 8316 50076
rect 8252 50016 8316 50020
rect 2352 49532 2416 49536
rect 2352 49476 2356 49532
rect 2356 49476 2412 49532
rect 2412 49476 2416 49532
rect 2352 49472 2416 49476
rect 2432 49532 2496 49536
rect 2432 49476 2436 49532
rect 2436 49476 2492 49532
rect 2492 49476 2496 49532
rect 2432 49472 2496 49476
rect 2512 49532 2576 49536
rect 2512 49476 2516 49532
rect 2516 49476 2572 49532
rect 2572 49476 2576 49532
rect 2512 49472 2576 49476
rect 2592 49532 2656 49536
rect 2592 49476 2596 49532
rect 2596 49476 2652 49532
rect 2652 49476 2656 49532
rect 2592 49472 2656 49476
rect 7352 49532 7416 49536
rect 7352 49476 7356 49532
rect 7356 49476 7412 49532
rect 7412 49476 7416 49532
rect 7352 49472 7416 49476
rect 7432 49532 7496 49536
rect 7432 49476 7436 49532
rect 7436 49476 7492 49532
rect 7492 49476 7496 49532
rect 7432 49472 7496 49476
rect 7512 49532 7576 49536
rect 7512 49476 7516 49532
rect 7516 49476 7572 49532
rect 7572 49476 7576 49532
rect 7512 49472 7576 49476
rect 7592 49532 7656 49536
rect 7592 49476 7596 49532
rect 7596 49476 7652 49532
rect 7652 49476 7656 49532
rect 7592 49472 7656 49476
rect 3012 48988 3076 48992
rect 3012 48932 3016 48988
rect 3016 48932 3072 48988
rect 3072 48932 3076 48988
rect 3012 48928 3076 48932
rect 3092 48988 3156 48992
rect 3092 48932 3096 48988
rect 3096 48932 3152 48988
rect 3152 48932 3156 48988
rect 3092 48928 3156 48932
rect 3172 48988 3236 48992
rect 3172 48932 3176 48988
rect 3176 48932 3232 48988
rect 3232 48932 3236 48988
rect 3172 48928 3236 48932
rect 3252 48988 3316 48992
rect 3252 48932 3256 48988
rect 3256 48932 3312 48988
rect 3312 48932 3316 48988
rect 3252 48928 3316 48932
rect 8012 48988 8076 48992
rect 8012 48932 8016 48988
rect 8016 48932 8072 48988
rect 8072 48932 8076 48988
rect 8012 48928 8076 48932
rect 8092 48988 8156 48992
rect 8092 48932 8096 48988
rect 8096 48932 8152 48988
rect 8152 48932 8156 48988
rect 8092 48928 8156 48932
rect 8172 48988 8236 48992
rect 8172 48932 8176 48988
rect 8176 48932 8232 48988
rect 8232 48932 8236 48988
rect 8172 48928 8236 48932
rect 8252 48988 8316 48992
rect 8252 48932 8256 48988
rect 8256 48932 8312 48988
rect 8312 48932 8316 48988
rect 8252 48928 8316 48932
rect 2352 48444 2416 48448
rect 2352 48388 2356 48444
rect 2356 48388 2412 48444
rect 2412 48388 2416 48444
rect 2352 48384 2416 48388
rect 2432 48444 2496 48448
rect 2432 48388 2436 48444
rect 2436 48388 2492 48444
rect 2492 48388 2496 48444
rect 2432 48384 2496 48388
rect 2512 48444 2576 48448
rect 2512 48388 2516 48444
rect 2516 48388 2572 48444
rect 2572 48388 2576 48444
rect 2512 48384 2576 48388
rect 2592 48444 2656 48448
rect 2592 48388 2596 48444
rect 2596 48388 2652 48444
rect 2652 48388 2656 48444
rect 2592 48384 2656 48388
rect 7352 48444 7416 48448
rect 7352 48388 7356 48444
rect 7356 48388 7412 48444
rect 7412 48388 7416 48444
rect 7352 48384 7416 48388
rect 7432 48444 7496 48448
rect 7432 48388 7436 48444
rect 7436 48388 7492 48444
rect 7492 48388 7496 48444
rect 7432 48384 7496 48388
rect 7512 48444 7576 48448
rect 7512 48388 7516 48444
rect 7516 48388 7572 48444
rect 7572 48388 7576 48444
rect 7512 48384 7576 48388
rect 7592 48444 7656 48448
rect 7592 48388 7596 48444
rect 7596 48388 7652 48444
rect 7652 48388 7656 48444
rect 7592 48384 7656 48388
rect 3012 47900 3076 47904
rect 3012 47844 3016 47900
rect 3016 47844 3072 47900
rect 3072 47844 3076 47900
rect 3012 47840 3076 47844
rect 3092 47900 3156 47904
rect 3092 47844 3096 47900
rect 3096 47844 3152 47900
rect 3152 47844 3156 47900
rect 3092 47840 3156 47844
rect 3172 47900 3236 47904
rect 3172 47844 3176 47900
rect 3176 47844 3232 47900
rect 3232 47844 3236 47900
rect 3172 47840 3236 47844
rect 3252 47900 3316 47904
rect 3252 47844 3256 47900
rect 3256 47844 3312 47900
rect 3312 47844 3316 47900
rect 3252 47840 3316 47844
rect 8012 47900 8076 47904
rect 8012 47844 8016 47900
rect 8016 47844 8072 47900
rect 8072 47844 8076 47900
rect 8012 47840 8076 47844
rect 8092 47900 8156 47904
rect 8092 47844 8096 47900
rect 8096 47844 8152 47900
rect 8152 47844 8156 47900
rect 8092 47840 8156 47844
rect 8172 47900 8236 47904
rect 8172 47844 8176 47900
rect 8176 47844 8232 47900
rect 8232 47844 8236 47900
rect 8172 47840 8236 47844
rect 8252 47900 8316 47904
rect 8252 47844 8256 47900
rect 8256 47844 8312 47900
rect 8312 47844 8316 47900
rect 8252 47840 8316 47844
rect 2352 47356 2416 47360
rect 2352 47300 2356 47356
rect 2356 47300 2412 47356
rect 2412 47300 2416 47356
rect 2352 47296 2416 47300
rect 2432 47356 2496 47360
rect 2432 47300 2436 47356
rect 2436 47300 2492 47356
rect 2492 47300 2496 47356
rect 2432 47296 2496 47300
rect 2512 47356 2576 47360
rect 2512 47300 2516 47356
rect 2516 47300 2572 47356
rect 2572 47300 2576 47356
rect 2512 47296 2576 47300
rect 2592 47356 2656 47360
rect 2592 47300 2596 47356
rect 2596 47300 2652 47356
rect 2652 47300 2656 47356
rect 2592 47296 2656 47300
rect 7352 47356 7416 47360
rect 7352 47300 7356 47356
rect 7356 47300 7412 47356
rect 7412 47300 7416 47356
rect 7352 47296 7416 47300
rect 7432 47356 7496 47360
rect 7432 47300 7436 47356
rect 7436 47300 7492 47356
rect 7492 47300 7496 47356
rect 7432 47296 7496 47300
rect 7512 47356 7576 47360
rect 7512 47300 7516 47356
rect 7516 47300 7572 47356
rect 7572 47300 7576 47356
rect 7512 47296 7576 47300
rect 7592 47356 7656 47360
rect 7592 47300 7596 47356
rect 7596 47300 7652 47356
rect 7652 47300 7656 47356
rect 7592 47296 7656 47300
rect 3012 46812 3076 46816
rect 3012 46756 3016 46812
rect 3016 46756 3072 46812
rect 3072 46756 3076 46812
rect 3012 46752 3076 46756
rect 3092 46812 3156 46816
rect 3092 46756 3096 46812
rect 3096 46756 3152 46812
rect 3152 46756 3156 46812
rect 3092 46752 3156 46756
rect 3172 46812 3236 46816
rect 3172 46756 3176 46812
rect 3176 46756 3232 46812
rect 3232 46756 3236 46812
rect 3172 46752 3236 46756
rect 3252 46812 3316 46816
rect 3252 46756 3256 46812
rect 3256 46756 3312 46812
rect 3312 46756 3316 46812
rect 3252 46752 3316 46756
rect 8012 46812 8076 46816
rect 8012 46756 8016 46812
rect 8016 46756 8072 46812
rect 8072 46756 8076 46812
rect 8012 46752 8076 46756
rect 8092 46812 8156 46816
rect 8092 46756 8096 46812
rect 8096 46756 8152 46812
rect 8152 46756 8156 46812
rect 8092 46752 8156 46756
rect 8172 46812 8236 46816
rect 8172 46756 8176 46812
rect 8176 46756 8232 46812
rect 8232 46756 8236 46812
rect 8172 46752 8236 46756
rect 8252 46812 8316 46816
rect 8252 46756 8256 46812
rect 8256 46756 8312 46812
rect 8312 46756 8316 46812
rect 8252 46752 8316 46756
rect 2352 46268 2416 46272
rect 2352 46212 2356 46268
rect 2356 46212 2412 46268
rect 2412 46212 2416 46268
rect 2352 46208 2416 46212
rect 2432 46268 2496 46272
rect 2432 46212 2436 46268
rect 2436 46212 2492 46268
rect 2492 46212 2496 46268
rect 2432 46208 2496 46212
rect 2512 46268 2576 46272
rect 2512 46212 2516 46268
rect 2516 46212 2572 46268
rect 2572 46212 2576 46268
rect 2512 46208 2576 46212
rect 2592 46268 2656 46272
rect 2592 46212 2596 46268
rect 2596 46212 2652 46268
rect 2652 46212 2656 46268
rect 2592 46208 2656 46212
rect 7352 46268 7416 46272
rect 7352 46212 7356 46268
rect 7356 46212 7412 46268
rect 7412 46212 7416 46268
rect 7352 46208 7416 46212
rect 7432 46268 7496 46272
rect 7432 46212 7436 46268
rect 7436 46212 7492 46268
rect 7492 46212 7496 46268
rect 7432 46208 7496 46212
rect 7512 46268 7576 46272
rect 7512 46212 7516 46268
rect 7516 46212 7572 46268
rect 7572 46212 7576 46268
rect 7512 46208 7576 46212
rect 7592 46268 7656 46272
rect 7592 46212 7596 46268
rect 7596 46212 7652 46268
rect 7652 46212 7656 46268
rect 7592 46208 7656 46212
rect 3012 45724 3076 45728
rect 3012 45668 3016 45724
rect 3016 45668 3072 45724
rect 3072 45668 3076 45724
rect 3012 45664 3076 45668
rect 3092 45724 3156 45728
rect 3092 45668 3096 45724
rect 3096 45668 3152 45724
rect 3152 45668 3156 45724
rect 3092 45664 3156 45668
rect 3172 45724 3236 45728
rect 3172 45668 3176 45724
rect 3176 45668 3232 45724
rect 3232 45668 3236 45724
rect 3172 45664 3236 45668
rect 3252 45724 3316 45728
rect 3252 45668 3256 45724
rect 3256 45668 3312 45724
rect 3312 45668 3316 45724
rect 3252 45664 3316 45668
rect 8012 45724 8076 45728
rect 8012 45668 8016 45724
rect 8016 45668 8072 45724
rect 8072 45668 8076 45724
rect 8012 45664 8076 45668
rect 8092 45724 8156 45728
rect 8092 45668 8096 45724
rect 8096 45668 8152 45724
rect 8152 45668 8156 45724
rect 8092 45664 8156 45668
rect 8172 45724 8236 45728
rect 8172 45668 8176 45724
rect 8176 45668 8232 45724
rect 8232 45668 8236 45724
rect 8172 45664 8236 45668
rect 8252 45724 8316 45728
rect 8252 45668 8256 45724
rect 8256 45668 8312 45724
rect 8312 45668 8316 45724
rect 8252 45664 8316 45668
rect 2352 45180 2416 45184
rect 2352 45124 2356 45180
rect 2356 45124 2412 45180
rect 2412 45124 2416 45180
rect 2352 45120 2416 45124
rect 2432 45180 2496 45184
rect 2432 45124 2436 45180
rect 2436 45124 2492 45180
rect 2492 45124 2496 45180
rect 2432 45120 2496 45124
rect 2512 45180 2576 45184
rect 2512 45124 2516 45180
rect 2516 45124 2572 45180
rect 2572 45124 2576 45180
rect 2512 45120 2576 45124
rect 2592 45180 2656 45184
rect 2592 45124 2596 45180
rect 2596 45124 2652 45180
rect 2652 45124 2656 45180
rect 2592 45120 2656 45124
rect 7352 45180 7416 45184
rect 7352 45124 7356 45180
rect 7356 45124 7412 45180
rect 7412 45124 7416 45180
rect 7352 45120 7416 45124
rect 7432 45180 7496 45184
rect 7432 45124 7436 45180
rect 7436 45124 7492 45180
rect 7492 45124 7496 45180
rect 7432 45120 7496 45124
rect 7512 45180 7576 45184
rect 7512 45124 7516 45180
rect 7516 45124 7572 45180
rect 7572 45124 7576 45180
rect 7512 45120 7576 45124
rect 7592 45180 7656 45184
rect 7592 45124 7596 45180
rect 7596 45124 7652 45180
rect 7652 45124 7656 45180
rect 7592 45120 7656 45124
rect 3012 44636 3076 44640
rect 3012 44580 3016 44636
rect 3016 44580 3072 44636
rect 3072 44580 3076 44636
rect 3012 44576 3076 44580
rect 3092 44636 3156 44640
rect 3092 44580 3096 44636
rect 3096 44580 3152 44636
rect 3152 44580 3156 44636
rect 3092 44576 3156 44580
rect 3172 44636 3236 44640
rect 3172 44580 3176 44636
rect 3176 44580 3232 44636
rect 3232 44580 3236 44636
rect 3172 44576 3236 44580
rect 3252 44636 3316 44640
rect 3252 44580 3256 44636
rect 3256 44580 3312 44636
rect 3312 44580 3316 44636
rect 3252 44576 3316 44580
rect 8012 44636 8076 44640
rect 8012 44580 8016 44636
rect 8016 44580 8072 44636
rect 8072 44580 8076 44636
rect 8012 44576 8076 44580
rect 8092 44636 8156 44640
rect 8092 44580 8096 44636
rect 8096 44580 8152 44636
rect 8152 44580 8156 44636
rect 8092 44576 8156 44580
rect 8172 44636 8236 44640
rect 8172 44580 8176 44636
rect 8176 44580 8232 44636
rect 8232 44580 8236 44636
rect 8172 44576 8236 44580
rect 8252 44636 8316 44640
rect 8252 44580 8256 44636
rect 8256 44580 8312 44636
rect 8312 44580 8316 44636
rect 8252 44576 8316 44580
rect 2352 44092 2416 44096
rect 2352 44036 2356 44092
rect 2356 44036 2412 44092
rect 2412 44036 2416 44092
rect 2352 44032 2416 44036
rect 2432 44092 2496 44096
rect 2432 44036 2436 44092
rect 2436 44036 2492 44092
rect 2492 44036 2496 44092
rect 2432 44032 2496 44036
rect 2512 44092 2576 44096
rect 2512 44036 2516 44092
rect 2516 44036 2572 44092
rect 2572 44036 2576 44092
rect 2512 44032 2576 44036
rect 2592 44092 2656 44096
rect 2592 44036 2596 44092
rect 2596 44036 2652 44092
rect 2652 44036 2656 44092
rect 2592 44032 2656 44036
rect 7352 44092 7416 44096
rect 7352 44036 7356 44092
rect 7356 44036 7412 44092
rect 7412 44036 7416 44092
rect 7352 44032 7416 44036
rect 7432 44092 7496 44096
rect 7432 44036 7436 44092
rect 7436 44036 7492 44092
rect 7492 44036 7496 44092
rect 7432 44032 7496 44036
rect 7512 44092 7576 44096
rect 7512 44036 7516 44092
rect 7516 44036 7572 44092
rect 7572 44036 7576 44092
rect 7512 44032 7576 44036
rect 7592 44092 7656 44096
rect 7592 44036 7596 44092
rect 7596 44036 7652 44092
rect 7652 44036 7656 44092
rect 7592 44032 7656 44036
rect 3012 43548 3076 43552
rect 3012 43492 3016 43548
rect 3016 43492 3072 43548
rect 3072 43492 3076 43548
rect 3012 43488 3076 43492
rect 3092 43548 3156 43552
rect 3092 43492 3096 43548
rect 3096 43492 3152 43548
rect 3152 43492 3156 43548
rect 3092 43488 3156 43492
rect 3172 43548 3236 43552
rect 3172 43492 3176 43548
rect 3176 43492 3232 43548
rect 3232 43492 3236 43548
rect 3172 43488 3236 43492
rect 3252 43548 3316 43552
rect 3252 43492 3256 43548
rect 3256 43492 3312 43548
rect 3312 43492 3316 43548
rect 3252 43488 3316 43492
rect 8012 43548 8076 43552
rect 8012 43492 8016 43548
rect 8016 43492 8072 43548
rect 8072 43492 8076 43548
rect 8012 43488 8076 43492
rect 8092 43548 8156 43552
rect 8092 43492 8096 43548
rect 8096 43492 8152 43548
rect 8152 43492 8156 43548
rect 8092 43488 8156 43492
rect 8172 43548 8236 43552
rect 8172 43492 8176 43548
rect 8176 43492 8232 43548
rect 8232 43492 8236 43548
rect 8172 43488 8236 43492
rect 8252 43548 8316 43552
rect 8252 43492 8256 43548
rect 8256 43492 8312 43548
rect 8312 43492 8316 43548
rect 8252 43488 8316 43492
rect 2352 43004 2416 43008
rect 2352 42948 2356 43004
rect 2356 42948 2412 43004
rect 2412 42948 2416 43004
rect 2352 42944 2416 42948
rect 2432 43004 2496 43008
rect 2432 42948 2436 43004
rect 2436 42948 2492 43004
rect 2492 42948 2496 43004
rect 2432 42944 2496 42948
rect 2512 43004 2576 43008
rect 2512 42948 2516 43004
rect 2516 42948 2572 43004
rect 2572 42948 2576 43004
rect 2512 42944 2576 42948
rect 2592 43004 2656 43008
rect 2592 42948 2596 43004
rect 2596 42948 2652 43004
rect 2652 42948 2656 43004
rect 2592 42944 2656 42948
rect 7352 43004 7416 43008
rect 7352 42948 7356 43004
rect 7356 42948 7412 43004
rect 7412 42948 7416 43004
rect 7352 42944 7416 42948
rect 7432 43004 7496 43008
rect 7432 42948 7436 43004
rect 7436 42948 7492 43004
rect 7492 42948 7496 43004
rect 7432 42944 7496 42948
rect 7512 43004 7576 43008
rect 7512 42948 7516 43004
rect 7516 42948 7572 43004
rect 7572 42948 7576 43004
rect 7512 42944 7576 42948
rect 7592 43004 7656 43008
rect 7592 42948 7596 43004
rect 7596 42948 7652 43004
rect 7652 42948 7656 43004
rect 7592 42944 7656 42948
rect 3012 42460 3076 42464
rect 3012 42404 3016 42460
rect 3016 42404 3072 42460
rect 3072 42404 3076 42460
rect 3012 42400 3076 42404
rect 3092 42460 3156 42464
rect 3092 42404 3096 42460
rect 3096 42404 3152 42460
rect 3152 42404 3156 42460
rect 3092 42400 3156 42404
rect 3172 42460 3236 42464
rect 3172 42404 3176 42460
rect 3176 42404 3232 42460
rect 3232 42404 3236 42460
rect 3172 42400 3236 42404
rect 3252 42460 3316 42464
rect 3252 42404 3256 42460
rect 3256 42404 3312 42460
rect 3312 42404 3316 42460
rect 3252 42400 3316 42404
rect 8012 42460 8076 42464
rect 8012 42404 8016 42460
rect 8016 42404 8072 42460
rect 8072 42404 8076 42460
rect 8012 42400 8076 42404
rect 8092 42460 8156 42464
rect 8092 42404 8096 42460
rect 8096 42404 8152 42460
rect 8152 42404 8156 42460
rect 8092 42400 8156 42404
rect 8172 42460 8236 42464
rect 8172 42404 8176 42460
rect 8176 42404 8232 42460
rect 8232 42404 8236 42460
rect 8172 42400 8236 42404
rect 8252 42460 8316 42464
rect 8252 42404 8256 42460
rect 8256 42404 8312 42460
rect 8312 42404 8316 42460
rect 8252 42400 8316 42404
rect 2352 41916 2416 41920
rect 2352 41860 2356 41916
rect 2356 41860 2412 41916
rect 2412 41860 2416 41916
rect 2352 41856 2416 41860
rect 2432 41916 2496 41920
rect 2432 41860 2436 41916
rect 2436 41860 2492 41916
rect 2492 41860 2496 41916
rect 2432 41856 2496 41860
rect 2512 41916 2576 41920
rect 2512 41860 2516 41916
rect 2516 41860 2572 41916
rect 2572 41860 2576 41916
rect 2512 41856 2576 41860
rect 2592 41916 2656 41920
rect 2592 41860 2596 41916
rect 2596 41860 2652 41916
rect 2652 41860 2656 41916
rect 2592 41856 2656 41860
rect 7352 41916 7416 41920
rect 7352 41860 7356 41916
rect 7356 41860 7412 41916
rect 7412 41860 7416 41916
rect 7352 41856 7416 41860
rect 7432 41916 7496 41920
rect 7432 41860 7436 41916
rect 7436 41860 7492 41916
rect 7492 41860 7496 41916
rect 7432 41856 7496 41860
rect 7512 41916 7576 41920
rect 7512 41860 7516 41916
rect 7516 41860 7572 41916
rect 7572 41860 7576 41916
rect 7512 41856 7576 41860
rect 7592 41916 7656 41920
rect 7592 41860 7596 41916
rect 7596 41860 7652 41916
rect 7652 41860 7656 41916
rect 7592 41856 7656 41860
rect 6316 41380 6380 41444
rect 3012 41372 3076 41376
rect 3012 41316 3016 41372
rect 3016 41316 3072 41372
rect 3072 41316 3076 41372
rect 3012 41312 3076 41316
rect 3092 41372 3156 41376
rect 3092 41316 3096 41372
rect 3096 41316 3152 41372
rect 3152 41316 3156 41372
rect 3092 41312 3156 41316
rect 3172 41372 3236 41376
rect 3172 41316 3176 41372
rect 3176 41316 3232 41372
rect 3232 41316 3236 41372
rect 3172 41312 3236 41316
rect 3252 41372 3316 41376
rect 3252 41316 3256 41372
rect 3256 41316 3312 41372
rect 3312 41316 3316 41372
rect 3252 41312 3316 41316
rect 8012 41372 8076 41376
rect 8012 41316 8016 41372
rect 8016 41316 8072 41372
rect 8072 41316 8076 41372
rect 8012 41312 8076 41316
rect 8092 41372 8156 41376
rect 8092 41316 8096 41372
rect 8096 41316 8152 41372
rect 8152 41316 8156 41372
rect 8092 41312 8156 41316
rect 8172 41372 8236 41376
rect 8172 41316 8176 41372
rect 8176 41316 8232 41372
rect 8232 41316 8236 41372
rect 8172 41312 8236 41316
rect 8252 41372 8316 41376
rect 8252 41316 8256 41372
rect 8256 41316 8312 41372
rect 8312 41316 8316 41372
rect 8252 41312 8316 41316
rect 2352 40828 2416 40832
rect 2352 40772 2356 40828
rect 2356 40772 2412 40828
rect 2412 40772 2416 40828
rect 2352 40768 2416 40772
rect 2432 40828 2496 40832
rect 2432 40772 2436 40828
rect 2436 40772 2492 40828
rect 2492 40772 2496 40828
rect 2432 40768 2496 40772
rect 2512 40828 2576 40832
rect 2512 40772 2516 40828
rect 2516 40772 2572 40828
rect 2572 40772 2576 40828
rect 2512 40768 2576 40772
rect 2592 40828 2656 40832
rect 2592 40772 2596 40828
rect 2596 40772 2652 40828
rect 2652 40772 2656 40828
rect 2592 40768 2656 40772
rect 7352 40828 7416 40832
rect 7352 40772 7356 40828
rect 7356 40772 7412 40828
rect 7412 40772 7416 40828
rect 7352 40768 7416 40772
rect 7432 40828 7496 40832
rect 7432 40772 7436 40828
rect 7436 40772 7492 40828
rect 7492 40772 7496 40828
rect 7432 40768 7496 40772
rect 7512 40828 7576 40832
rect 7512 40772 7516 40828
rect 7516 40772 7572 40828
rect 7572 40772 7576 40828
rect 7512 40768 7576 40772
rect 7592 40828 7656 40832
rect 7592 40772 7596 40828
rect 7596 40772 7652 40828
rect 7652 40772 7656 40828
rect 7592 40768 7656 40772
rect 3012 40284 3076 40288
rect 3012 40228 3016 40284
rect 3016 40228 3072 40284
rect 3072 40228 3076 40284
rect 3012 40224 3076 40228
rect 3092 40284 3156 40288
rect 3092 40228 3096 40284
rect 3096 40228 3152 40284
rect 3152 40228 3156 40284
rect 3092 40224 3156 40228
rect 3172 40284 3236 40288
rect 3172 40228 3176 40284
rect 3176 40228 3232 40284
rect 3232 40228 3236 40284
rect 3172 40224 3236 40228
rect 3252 40284 3316 40288
rect 3252 40228 3256 40284
rect 3256 40228 3312 40284
rect 3312 40228 3316 40284
rect 3252 40224 3316 40228
rect 8012 40284 8076 40288
rect 8012 40228 8016 40284
rect 8016 40228 8072 40284
rect 8072 40228 8076 40284
rect 8012 40224 8076 40228
rect 8092 40284 8156 40288
rect 8092 40228 8096 40284
rect 8096 40228 8152 40284
rect 8152 40228 8156 40284
rect 8092 40224 8156 40228
rect 8172 40284 8236 40288
rect 8172 40228 8176 40284
rect 8176 40228 8232 40284
rect 8232 40228 8236 40284
rect 8172 40224 8236 40228
rect 8252 40284 8316 40288
rect 8252 40228 8256 40284
rect 8256 40228 8312 40284
rect 8312 40228 8316 40284
rect 8252 40224 8316 40228
rect 6684 40020 6748 40084
rect 2352 39740 2416 39744
rect 2352 39684 2356 39740
rect 2356 39684 2412 39740
rect 2412 39684 2416 39740
rect 2352 39680 2416 39684
rect 2432 39740 2496 39744
rect 2432 39684 2436 39740
rect 2436 39684 2492 39740
rect 2492 39684 2496 39740
rect 2432 39680 2496 39684
rect 2512 39740 2576 39744
rect 2512 39684 2516 39740
rect 2516 39684 2572 39740
rect 2572 39684 2576 39740
rect 2512 39680 2576 39684
rect 2592 39740 2656 39744
rect 2592 39684 2596 39740
rect 2596 39684 2652 39740
rect 2652 39684 2656 39740
rect 2592 39680 2656 39684
rect 7352 39740 7416 39744
rect 7352 39684 7356 39740
rect 7356 39684 7412 39740
rect 7412 39684 7416 39740
rect 7352 39680 7416 39684
rect 7432 39740 7496 39744
rect 7432 39684 7436 39740
rect 7436 39684 7492 39740
rect 7492 39684 7496 39740
rect 7432 39680 7496 39684
rect 7512 39740 7576 39744
rect 7512 39684 7516 39740
rect 7516 39684 7572 39740
rect 7572 39684 7576 39740
rect 7512 39680 7576 39684
rect 7592 39740 7656 39744
rect 7592 39684 7596 39740
rect 7596 39684 7652 39740
rect 7652 39684 7656 39740
rect 7592 39680 7656 39684
rect 3012 39196 3076 39200
rect 3012 39140 3016 39196
rect 3016 39140 3072 39196
rect 3072 39140 3076 39196
rect 3012 39136 3076 39140
rect 3092 39196 3156 39200
rect 3092 39140 3096 39196
rect 3096 39140 3152 39196
rect 3152 39140 3156 39196
rect 3092 39136 3156 39140
rect 3172 39196 3236 39200
rect 3172 39140 3176 39196
rect 3176 39140 3232 39196
rect 3232 39140 3236 39196
rect 3172 39136 3236 39140
rect 3252 39196 3316 39200
rect 3252 39140 3256 39196
rect 3256 39140 3312 39196
rect 3312 39140 3316 39196
rect 3252 39136 3316 39140
rect 8012 39196 8076 39200
rect 8012 39140 8016 39196
rect 8016 39140 8072 39196
rect 8072 39140 8076 39196
rect 8012 39136 8076 39140
rect 8092 39196 8156 39200
rect 8092 39140 8096 39196
rect 8096 39140 8152 39196
rect 8152 39140 8156 39196
rect 8092 39136 8156 39140
rect 8172 39196 8236 39200
rect 8172 39140 8176 39196
rect 8176 39140 8232 39196
rect 8232 39140 8236 39196
rect 8172 39136 8236 39140
rect 8252 39196 8316 39200
rect 8252 39140 8256 39196
rect 8256 39140 8312 39196
rect 8312 39140 8316 39196
rect 8252 39136 8316 39140
rect 2352 38652 2416 38656
rect 2352 38596 2356 38652
rect 2356 38596 2412 38652
rect 2412 38596 2416 38652
rect 2352 38592 2416 38596
rect 2432 38652 2496 38656
rect 2432 38596 2436 38652
rect 2436 38596 2492 38652
rect 2492 38596 2496 38652
rect 2432 38592 2496 38596
rect 2512 38652 2576 38656
rect 2512 38596 2516 38652
rect 2516 38596 2572 38652
rect 2572 38596 2576 38652
rect 2512 38592 2576 38596
rect 2592 38652 2656 38656
rect 2592 38596 2596 38652
rect 2596 38596 2652 38652
rect 2652 38596 2656 38652
rect 2592 38592 2656 38596
rect 7352 38652 7416 38656
rect 7352 38596 7356 38652
rect 7356 38596 7412 38652
rect 7412 38596 7416 38652
rect 7352 38592 7416 38596
rect 7432 38652 7496 38656
rect 7432 38596 7436 38652
rect 7436 38596 7492 38652
rect 7492 38596 7496 38652
rect 7432 38592 7496 38596
rect 7512 38652 7576 38656
rect 7512 38596 7516 38652
rect 7516 38596 7572 38652
rect 7572 38596 7576 38652
rect 7512 38592 7576 38596
rect 7592 38652 7656 38656
rect 7592 38596 7596 38652
rect 7596 38596 7652 38652
rect 7652 38596 7656 38652
rect 7592 38592 7656 38596
rect 3012 38108 3076 38112
rect 3012 38052 3016 38108
rect 3016 38052 3072 38108
rect 3072 38052 3076 38108
rect 3012 38048 3076 38052
rect 3092 38108 3156 38112
rect 3092 38052 3096 38108
rect 3096 38052 3152 38108
rect 3152 38052 3156 38108
rect 3092 38048 3156 38052
rect 3172 38108 3236 38112
rect 3172 38052 3176 38108
rect 3176 38052 3232 38108
rect 3232 38052 3236 38108
rect 3172 38048 3236 38052
rect 3252 38108 3316 38112
rect 3252 38052 3256 38108
rect 3256 38052 3312 38108
rect 3312 38052 3316 38108
rect 3252 38048 3316 38052
rect 8012 38108 8076 38112
rect 8012 38052 8016 38108
rect 8016 38052 8072 38108
rect 8072 38052 8076 38108
rect 8012 38048 8076 38052
rect 8092 38108 8156 38112
rect 8092 38052 8096 38108
rect 8096 38052 8152 38108
rect 8152 38052 8156 38108
rect 8092 38048 8156 38052
rect 8172 38108 8236 38112
rect 8172 38052 8176 38108
rect 8176 38052 8232 38108
rect 8232 38052 8236 38108
rect 8172 38048 8236 38052
rect 8252 38108 8316 38112
rect 8252 38052 8256 38108
rect 8256 38052 8312 38108
rect 8312 38052 8316 38108
rect 8252 38048 8316 38052
rect 2352 37564 2416 37568
rect 2352 37508 2356 37564
rect 2356 37508 2412 37564
rect 2412 37508 2416 37564
rect 2352 37504 2416 37508
rect 2432 37564 2496 37568
rect 2432 37508 2436 37564
rect 2436 37508 2492 37564
rect 2492 37508 2496 37564
rect 2432 37504 2496 37508
rect 2512 37564 2576 37568
rect 2512 37508 2516 37564
rect 2516 37508 2572 37564
rect 2572 37508 2576 37564
rect 2512 37504 2576 37508
rect 2592 37564 2656 37568
rect 2592 37508 2596 37564
rect 2596 37508 2652 37564
rect 2652 37508 2656 37564
rect 2592 37504 2656 37508
rect 7352 37564 7416 37568
rect 7352 37508 7356 37564
rect 7356 37508 7412 37564
rect 7412 37508 7416 37564
rect 7352 37504 7416 37508
rect 7432 37564 7496 37568
rect 7432 37508 7436 37564
rect 7436 37508 7492 37564
rect 7492 37508 7496 37564
rect 7432 37504 7496 37508
rect 7512 37564 7576 37568
rect 7512 37508 7516 37564
rect 7516 37508 7572 37564
rect 7572 37508 7576 37564
rect 7512 37504 7576 37508
rect 7592 37564 7656 37568
rect 7592 37508 7596 37564
rect 7596 37508 7652 37564
rect 7652 37508 7656 37564
rect 7592 37504 7656 37508
rect 3012 37020 3076 37024
rect 3012 36964 3016 37020
rect 3016 36964 3072 37020
rect 3072 36964 3076 37020
rect 3012 36960 3076 36964
rect 3092 37020 3156 37024
rect 3092 36964 3096 37020
rect 3096 36964 3152 37020
rect 3152 36964 3156 37020
rect 3092 36960 3156 36964
rect 3172 37020 3236 37024
rect 3172 36964 3176 37020
rect 3176 36964 3232 37020
rect 3232 36964 3236 37020
rect 3172 36960 3236 36964
rect 3252 37020 3316 37024
rect 3252 36964 3256 37020
rect 3256 36964 3312 37020
rect 3312 36964 3316 37020
rect 3252 36960 3316 36964
rect 8012 37020 8076 37024
rect 8012 36964 8016 37020
rect 8016 36964 8072 37020
rect 8072 36964 8076 37020
rect 8012 36960 8076 36964
rect 8092 37020 8156 37024
rect 8092 36964 8096 37020
rect 8096 36964 8152 37020
rect 8152 36964 8156 37020
rect 8092 36960 8156 36964
rect 8172 37020 8236 37024
rect 8172 36964 8176 37020
rect 8176 36964 8232 37020
rect 8232 36964 8236 37020
rect 8172 36960 8236 36964
rect 8252 37020 8316 37024
rect 8252 36964 8256 37020
rect 8256 36964 8312 37020
rect 8312 36964 8316 37020
rect 8252 36960 8316 36964
rect 2352 36476 2416 36480
rect 2352 36420 2356 36476
rect 2356 36420 2412 36476
rect 2412 36420 2416 36476
rect 2352 36416 2416 36420
rect 2432 36476 2496 36480
rect 2432 36420 2436 36476
rect 2436 36420 2492 36476
rect 2492 36420 2496 36476
rect 2432 36416 2496 36420
rect 2512 36476 2576 36480
rect 2512 36420 2516 36476
rect 2516 36420 2572 36476
rect 2572 36420 2576 36476
rect 2512 36416 2576 36420
rect 2592 36476 2656 36480
rect 2592 36420 2596 36476
rect 2596 36420 2652 36476
rect 2652 36420 2656 36476
rect 2592 36416 2656 36420
rect 7352 36476 7416 36480
rect 7352 36420 7356 36476
rect 7356 36420 7412 36476
rect 7412 36420 7416 36476
rect 7352 36416 7416 36420
rect 7432 36476 7496 36480
rect 7432 36420 7436 36476
rect 7436 36420 7492 36476
rect 7492 36420 7496 36476
rect 7432 36416 7496 36420
rect 7512 36476 7576 36480
rect 7512 36420 7516 36476
rect 7516 36420 7572 36476
rect 7572 36420 7576 36476
rect 7512 36416 7576 36420
rect 7592 36476 7656 36480
rect 7592 36420 7596 36476
rect 7596 36420 7652 36476
rect 7652 36420 7656 36476
rect 7592 36416 7656 36420
rect 3012 35932 3076 35936
rect 3012 35876 3016 35932
rect 3016 35876 3072 35932
rect 3072 35876 3076 35932
rect 3012 35872 3076 35876
rect 3092 35932 3156 35936
rect 3092 35876 3096 35932
rect 3096 35876 3152 35932
rect 3152 35876 3156 35932
rect 3092 35872 3156 35876
rect 3172 35932 3236 35936
rect 3172 35876 3176 35932
rect 3176 35876 3232 35932
rect 3232 35876 3236 35932
rect 3172 35872 3236 35876
rect 3252 35932 3316 35936
rect 3252 35876 3256 35932
rect 3256 35876 3312 35932
rect 3312 35876 3316 35932
rect 3252 35872 3316 35876
rect 8012 35932 8076 35936
rect 8012 35876 8016 35932
rect 8016 35876 8072 35932
rect 8072 35876 8076 35932
rect 8012 35872 8076 35876
rect 8092 35932 8156 35936
rect 8092 35876 8096 35932
rect 8096 35876 8152 35932
rect 8152 35876 8156 35932
rect 8092 35872 8156 35876
rect 8172 35932 8236 35936
rect 8172 35876 8176 35932
rect 8176 35876 8232 35932
rect 8232 35876 8236 35932
rect 8172 35872 8236 35876
rect 8252 35932 8316 35936
rect 8252 35876 8256 35932
rect 8256 35876 8312 35932
rect 8312 35876 8316 35932
rect 8252 35872 8316 35876
rect 2352 35388 2416 35392
rect 2352 35332 2356 35388
rect 2356 35332 2412 35388
rect 2412 35332 2416 35388
rect 2352 35328 2416 35332
rect 2432 35388 2496 35392
rect 2432 35332 2436 35388
rect 2436 35332 2492 35388
rect 2492 35332 2496 35388
rect 2432 35328 2496 35332
rect 2512 35388 2576 35392
rect 2512 35332 2516 35388
rect 2516 35332 2572 35388
rect 2572 35332 2576 35388
rect 2512 35328 2576 35332
rect 2592 35388 2656 35392
rect 2592 35332 2596 35388
rect 2596 35332 2652 35388
rect 2652 35332 2656 35388
rect 2592 35328 2656 35332
rect 7352 35388 7416 35392
rect 7352 35332 7356 35388
rect 7356 35332 7412 35388
rect 7412 35332 7416 35388
rect 7352 35328 7416 35332
rect 7432 35388 7496 35392
rect 7432 35332 7436 35388
rect 7436 35332 7492 35388
rect 7492 35332 7496 35388
rect 7432 35328 7496 35332
rect 7512 35388 7576 35392
rect 7512 35332 7516 35388
rect 7516 35332 7572 35388
rect 7572 35332 7576 35388
rect 7512 35328 7576 35332
rect 7592 35388 7656 35392
rect 7592 35332 7596 35388
rect 7596 35332 7652 35388
rect 7652 35332 7656 35388
rect 7592 35328 7656 35332
rect 3012 34844 3076 34848
rect 3012 34788 3016 34844
rect 3016 34788 3072 34844
rect 3072 34788 3076 34844
rect 3012 34784 3076 34788
rect 3092 34844 3156 34848
rect 3092 34788 3096 34844
rect 3096 34788 3152 34844
rect 3152 34788 3156 34844
rect 3092 34784 3156 34788
rect 3172 34844 3236 34848
rect 3172 34788 3176 34844
rect 3176 34788 3232 34844
rect 3232 34788 3236 34844
rect 3172 34784 3236 34788
rect 3252 34844 3316 34848
rect 3252 34788 3256 34844
rect 3256 34788 3312 34844
rect 3312 34788 3316 34844
rect 3252 34784 3316 34788
rect 8012 34844 8076 34848
rect 8012 34788 8016 34844
rect 8016 34788 8072 34844
rect 8072 34788 8076 34844
rect 8012 34784 8076 34788
rect 8092 34844 8156 34848
rect 8092 34788 8096 34844
rect 8096 34788 8152 34844
rect 8152 34788 8156 34844
rect 8092 34784 8156 34788
rect 8172 34844 8236 34848
rect 8172 34788 8176 34844
rect 8176 34788 8232 34844
rect 8232 34788 8236 34844
rect 8172 34784 8236 34788
rect 8252 34844 8316 34848
rect 8252 34788 8256 34844
rect 8256 34788 8312 34844
rect 8312 34788 8316 34844
rect 8252 34784 8316 34788
rect 2352 34300 2416 34304
rect 2352 34244 2356 34300
rect 2356 34244 2412 34300
rect 2412 34244 2416 34300
rect 2352 34240 2416 34244
rect 2432 34300 2496 34304
rect 2432 34244 2436 34300
rect 2436 34244 2492 34300
rect 2492 34244 2496 34300
rect 2432 34240 2496 34244
rect 2512 34300 2576 34304
rect 2512 34244 2516 34300
rect 2516 34244 2572 34300
rect 2572 34244 2576 34300
rect 2512 34240 2576 34244
rect 2592 34300 2656 34304
rect 2592 34244 2596 34300
rect 2596 34244 2652 34300
rect 2652 34244 2656 34300
rect 2592 34240 2656 34244
rect 7352 34300 7416 34304
rect 7352 34244 7356 34300
rect 7356 34244 7412 34300
rect 7412 34244 7416 34300
rect 7352 34240 7416 34244
rect 7432 34300 7496 34304
rect 7432 34244 7436 34300
rect 7436 34244 7492 34300
rect 7492 34244 7496 34300
rect 7432 34240 7496 34244
rect 7512 34300 7576 34304
rect 7512 34244 7516 34300
rect 7516 34244 7572 34300
rect 7572 34244 7576 34300
rect 7512 34240 7576 34244
rect 7592 34300 7656 34304
rect 7592 34244 7596 34300
rect 7596 34244 7652 34300
rect 7652 34244 7656 34300
rect 7592 34240 7656 34244
rect 3012 33756 3076 33760
rect 3012 33700 3016 33756
rect 3016 33700 3072 33756
rect 3072 33700 3076 33756
rect 3012 33696 3076 33700
rect 3092 33756 3156 33760
rect 3092 33700 3096 33756
rect 3096 33700 3152 33756
rect 3152 33700 3156 33756
rect 3092 33696 3156 33700
rect 3172 33756 3236 33760
rect 3172 33700 3176 33756
rect 3176 33700 3232 33756
rect 3232 33700 3236 33756
rect 3172 33696 3236 33700
rect 3252 33756 3316 33760
rect 3252 33700 3256 33756
rect 3256 33700 3312 33756
rect 3312 33700 3316 33756
rect 3252 33696 3316 33700
rect 8012 33756 8076 33760
rect 8012 33700 8016 33756
rect 8016 33700 8072 33756
rect 8072 33700 8076 33756
rect 8012 33696 8076 33700
rect 8092 33756 8156 33760
rect 8092 33700 8096 33756
rect 8096 33700 8152 33756
rect 8152 33700 8156 33756
rect 8092 33696 8156 33700
rect 8172 33756 8236 33760
rect 8172 33700 8176 33756
rect 8176 33700 8232 33756
rect 8232 33700 8236 33756
rect 8172 33696 8236 33700
rect 8252 33756 8316 33760
rect 8252 33700 8256 33756
rect 8256 33700 8312 33756
rect 8312 33700 8316 33756
rect 8252 33696 8316 33700
rect 2352 33212 2416 33216
rect 2352 33156 2356 33212
rect 2356 33156 2412 33212
rect 2412 33156 2416 33212
rect 2352 33152 2416 33156
rect 2432 33212 2496 33216
rect 2432 33156 2436 33212
rect 2436 33156 2492 33212
rect 2492 33156 2496 33212
rect 2432 33152 2496 33156
rect 2512 33212 2576 33216
rect 2512 33156 2516 33212
rect 2516 33156 2572 33212
rect 2572 33156 2576 33212
rect 2512 33152 2576 33156
rect 2592 33212 2656 33216
rect 2592 33156 2596 33212
rect 2596 33156 2652 33212
rect 2652 33156 2656 33212
rect 2592 33152 2656 33156
rect 7352 33212 7416 33216
rect 7352 33156 7356 33212
rect 7356 33156 7412 33212
rect 7412 33156 7416 33212
rect 7352 33152 7416 33156
rect 7432 33212 7496 33216
rect 7432 33156 7436 33212
rect 7436 33156 7492 33212
rect 7492 33156 7496 33212
rect 7432 33152 7496 33156
rect 7512 33212 7576 33216
rect 7512 33156 7516 33212
rect 7516 33156 7572 33212
rect 7572 33156 7576 33212
rect 7512 33152 7576 33156
rect 7592 33212 7656 33216
rect 7592 33156 7596 33212
rect 7596 33156 7652 33212
rect 7652 33156 7656 33212
rect 7592 33152 7656 33156
rect 3012 32668 3076 32672
rect 3012 32612 3016 32668
rect 3016 32612 3072 32668
rect 3072 32612 3076 32668
rect 3012 32608 3076 32612
rect 3092 32668 3156 32672
rect 3092 32612 3096 32668
rect 3096 32612 3152 32668
rect 3152 32612 3156 32668
rect 3092 32608 3156 32612
rect 3172 32668 3236 32672
rect 3172 32612 3176 32668
rect 3176 32612 3232 32668
rect 3232 32612 3236 32668
rect 3172 32608 3236 32612
rect 3252 32668 3316 32672
rect 3252 32612 3256 32668
rect 3256 32612 3312 32668
rect 3312 32612 3316 32668
rect 3252 32608 3316 32612
rect 8012 32668 8076 32672
rect 8012 32612 8016 32668
rect 8016 32612 8072 32668
rect 8072 32612 8076 32668
rect 8012 32608 8076 32612
rect 8092 32668 8156 32672
rect 8092 32612 8096 32668
rect 8096 32612 8152 32668
rect 8152 32612 8156 32668
rect 8092 32608 8156 32612
rect 8172 32668 8236 32672
rect 8172 32612 8176 32668
rect 8176 32612 8232 32668
rect 8232 32612 8236 32668
rect 8172 32608 8236 32612
rect 8252 32668 8316 32672
rect 8252 32612 8256 32668
rect 8256 32612 8312 32668
rect 8312 32612 8316 32668
rect 8252 32608 8316 32612
rect 2352 32124 2416 32128
rect 2352 32068 2356 32124
rect 2356 32068 2412 32124
rect 2412 32068 2416 32124
rect 2352 32064 2416 32068
rect 2432 32124 2496 32128
rect 2432 32068 2436 32124
rect 2436 32068 2492 32124
rect 2492 32068 2496 32124
rect 2432 32064 2496 32068
rect 2512 32124 2576 32128
rect 2512 32068 2516 32124
rect 2516 32068 2572 32124
rect 2572 32068 2576 32124
rect 2512 32064 2576 32068
rect 2592 32124 2656 32128
rect 2592 32068 2596 32124
rect 2596 32068 2652 32124
rect 2652 32068 2656 32124
rect 2592 32064 2656 32068
rect 7352 32124 7416 32128
rect 7352 32068 7356 32124
rect 7356 32068 7412 32124
rect 7412 32068 7416 32124
rect 7352 32064 7416 32068
rect 7432 32124 7496 32128
rect 7432 32068 7436 32124
rect 7436 32068 7492 32124
rect 7492 32068 7496 32124
rect 7432 32064 7496 32068
rect 7512 32124 7576 32128
rect 7512 32068 7516 32124
rect 7516 32068 7572 32124
rect 7572 32068 7576 32124
rect 7512 32064 7576 32068
rect 7592 32124 7656 32128
rect 7592 32068 7596 32124
rect 7596 32068 7652 32124
rect 7652 32068 7656 32124
rect 7592 32064 7656 32068
rect 3012 31580 3076 31584
rect 3012 31524 3016 31580
rect 3016 31524 3072 31580
rect 3072 31524 3076 31580
rect 3012 31520 3076 31524
rect 3092 31580 3156 31584
rect 3092 31524 3096 31580
rect 3096 31524 3152 31580
rect 3152 31524 3156 31580
rect 3092 31520 3156 31524
rect 3172 31580 3236 31584
rect 3172 31524 3176 31580
rect 3176 31524 3232 31580
rect 3232 31524 3236 31580
rect 3172 31520 3236 31524
rect 3252 31580 3316 31584
rect 3252 31524 3256 31580
rect 3256 31524 3312 31580
rect 3312 31524 3316 31580
rect 3252 31520 3316 31524
rect 8012 31580 8076 31584
rect 8012 31524 8016 31580
rect 8016 31524 8072 31580
rect 8072 31524 8076 31580
rect 8012 31520 8076 31524
rect 8092 31580 8156 31584
rect 8092 31524 8096 31580
rect 8096 31524 8152 31580
rect 8152 31524 8156 31580
rect 8092 31520 8156 31524
rect 8172 31580 8236 31584
rect 8172 31524 8176 31580
rect 8176 31524 8232 31580
rect 8232 31524 8236 31580
rect 8172 31520 8236 31524
rect 8252 31580 8316 31584
rect 8252 31524 8256 31580
rect 8256 31524 8312 31580
rect 8312 31524 8316 31580
rect 8252 31520 8316 31524
rect 2352 31036 2416 31040
rect 2352 30980 2356 31036
rect 2356 30980 2412 31036
rect 2412 30980 2416 31036
rect 2352 30976 2416 30980
rect 2432 31036 2496 31040
rect 2432 30980 2436 31036
rect 2436 30980 2492 31036
rect 2492 30980 2496 31036
rect 2432 30976 2496 30980
rect 2512 31036 2576 31040
rect 2512 30980 2516 31036
rect 2516 30980 2572 31036
rect 2572 30980 2576 31036
rect 2512 30976 2576 30980
rect 2592 31036 2656 31040
rect 2592 30980 2596 31036
rect 2596 30980 2652 31036
rect 2652 30980 2656 31036
rect 2592 30976 2656 30980
rect 7352 31036 7416 31040
rect 7352 30980 7356 31036
rect 7356 30980 7412 31036
rect 7412 30980 7416 31036
rect 7352 30976 7416 30980
rect 7432 31036 7496 31040
rect 7432 30980 7436 31036
rect 7436 30980 7492 31036
rect 7492 30980 7496 31036
rect 7432 30976 7496 30980
rect 7512 31036 7576 31040
rect 7512 30980 7516 31036
rect 7516 30980 7572 31036
rect 7572 30980 7576 31036
rect 7512 30976 7576 30980
rect 7592 31036 7656 31040
rect 7592 30980 7596 31036
rect 7596 30980 7652 31036
rect 7652 30980 7656 31036
rect 7592 30976 7656 30980
rect 3012 30492 3076 30496
rect 3012 30436 3016 30492
rect 3016 30436 3072 30492
rect 3072 30436 3076 30492
rect 3012 30432 3076 30436
rect 3092 30492 3156 30496
rect 3092 30436 3096 30492
rect 3096 30436 3152 30492
rect 3152 30436 3156 30492
rect 3092 30432 3156 30436
rect 3172 30492 3236 30496
rect 3172 30436 3176 30492
rect 3176 30436 3232 30492
rect 3232 30436 3236 30492
rect 3172 30432 3236 30436
rect 3252 30492 3316 30496
rect 3252 30436 3256 30492
rect 3256 30436 3312 30492
rect 3312 30436 3316 30492
rect 3252 30432 3316 30436
rect 8012 30492 8076 30496
rect 8012 30436 8016 30492
rect 8016 30436 8072 30492
rect 8072 30436 8076 30492
rect 8012 30432 8076 30436
rect 8092 30492 8156 30496
rect 8092 30436 8096 30492
rect 8096 30436 8152 30492
rect 8152 30436 8156 30492
rect 8092 30432 8156 30436
rect 8172 30492 8236 30496
rect 8172 30436 8176 30492
rect 8176 30436 8232 30492
rect 8232 30436 8236 30492
rect 8172 30432 8236 30436
rect 8252 30492 8316 30496
rect 8252 30436 8256 30492
rect 8256 30436 8312 30492
rect 8312 30436 8316 30492
rect 8252 30432 8316 30436
rect 2352 29948 2416 29952
rect 2352 29892 2356 29948
rect 2356 29892 2412 29948
rect 2412 29892 2416 29948
rect 2352 29888 2416 29892
rect 2432 29948 2496 29952
rect 2432 29892 2436 29948
rect 2436 29892 2492 29948
rect 2492 29892 2496 29948
rect 2432 29888 2496 29892
rect 2512 29948 2576 29952
rect 2512 29892 2516 29948
rect 2516 29892 2572 29948
rect 2572 29892 2576 29948
rect 2512 29888 2576 29892
rect 2592 29948 2656 29952
rect 2592 29892 2596 29948
rect 2596 29892 2652 29948
rect 2652 29892 2656 29948
rect 2592 29888 2656 29892
rect 7352 29948 7416 29952
rect 7352 29892 7356 29948
rect 7356 29892 7412 29948
rect 7412 29892 7416 29948
rect 7352 29888 7416 29892
rect 7432 29948 7496 29952
rect 7432 29892 7436 29948
rect 7436 29892 7492 29948
rect 7492 29892 7496 29948
rect 7432 29888 7496 29892
rect 7512 29948 7576 29952
rect 7512 29892 7516 29948
rect 7516 29892 7572 29948
rect 7572 29892 7576 29948
rect 7512 29888 7576 29892
rect 7592 29948 7656 29952
rect 7592 29892 7596 29948
rect 7596 29892 7652 29948
rect 7652 29892 7656 29948
rect 7592 29888 7656 29892
rect 3012 29404 3076 29408
rect 3012 29348 3016 29404
rect 3016 29348 3072 29404
rect 3072 29348 3076 29404
rect 3012 29344 3076 29348
rect 3092 29404 3156 29408
rect 3092 29348 3096 29404
rect 3096 29348 3152 29404
rect 3152 29348 3156 29404
rect 3092 29344 3156 29348
rect 3172 29404 3236 29408
rect 3172 29348 3176 29404
rect 3176 29348 3232 29404
rect 3232 29348 3236 29404
rect 3172 29344 3236 29348
rect 3252 29404 3316 29408
rect 3252 29348 3256 29404
rect 3256 29348 3312 29404
rect 3312 29348 3316 29404
rect 3252 29344 3316 29348
rect 8012 29404 8076 29408
rect 8012 29348 8016 29404
rect 8016 29348 8072 29404
rect 8072 29348 8076 29404
rect 8012 29344 8076 29348
rect 8092 29404 8156 29408
rect 8092 29348 8096 29404
rect 8096 29348 8152 29404
rect 8152 29348 8156 29404
rect 8092 29344 8156 29348
rect 8172 29404 8236 29408
rect 8172 29348 8176 29404
rect 8176 29348 8232 29404
rect 8232 29348 8236 29404
rect 8172 29344 8236 29348
rect 8252 29404 8316 29408
rect 8252 29348 8256 29404
rect 8256 29348 8312 29404
rect 8312 29348 8316 29404
rect 8252 29344 8316 29348
rect 2352 28860 2416 28864
rect 2352 28804 2356 28860
rect 2356 28804 2412 28860
rect 2412 28804 2416 28860
rect 2352 28800 2416 28804
rect 2432 28860 2496 28864
rect 2432 28804 2436 28860
rect 2436 28804 2492 28860
rect 2492 28804 2496 28860
rect 2432 28800 2496 28804
rect 2512 28860 2576 28864
rect 2512 28804 2516 28860
rect 2516 28804 2572 28860
rect 2572 28804 2576 28860
rect 2512 28800 2576 28804
rect 2592 28860 2656 28864
rect 2592 28804 2596 28860
rect 2596 28804 2652 28860
rect 2652 28804 2656 28860
rect 2592 28800 2656 28804
rect 7352 28860 7416 28864
rect 7352 28804 7356 28860
rect 7356 28804 7412 28860
rect 7412 28804 7416 28860
rect 7352 28800 7416 28804
rect 7432 28860 7496 28864
rect 7432 28804 7436 28860
rect 7436 28804 7492 28860
rect 7492 28804 7496 28860
rect 7432 28800 7496 28804
rect 7512 28860 7576 28864
rect 7512 28804 7516 28860
rect 7516 28804 7572 28860
rect 7572 28804 7576 28860
rect 7512 28800 7576 28804
rect 7592 28860 7656 28864
rect 7592 28804 7596 28860
rect 7596 28804 7652 28860
rect 7652 28804 7656 28860
rect 7592 28800 7656 28804
rect 3012 28316 3076 28320
rect 3012 28260 3016 28316
rect 3016 28260 3072 28316
rect 3072 28260 3076 28316
rect 3012 28256 3076 28260
rect 3092 28316 3156 28320
rect 3092 28260 3096 28316
rect 3096 28260 3152 28316
rect 3152 28260 3156 28316
rect 3092 28256 3156 28260
rect 3172 28316 3236 28320
rect 3172 28260 3176 28316
rect 3176 28260 3232 28316
rect 3232 28260 3236 28316
rect 3172 28256 3236 28260
rect 3252 28316 3316 28320
rect 3252 28260 3256 28316
rect 3256 28260 3312 28316
rect 3312 28260 3316 28316
rect 3252 28256 3316 28260
rect 8012 28316 8076 28320
rect 8012 28260 8016 28316
rect 8016 28260 8072 28316
rect 8072 28260 8076 28316
rect 8012 28256 8076 28260
rect 8092 28316 8156 28320
rect 8092 28260 8096 28316
rect 8096 28260 8152 28316
rect 8152 28260 8156 28316
rect 8092 28256 8156 28260
rect 8172 28316 8236 28320
rect 8172 28260 8176 28316
rect 8176 28260 8232 28316
rect 8232 28260 8236 28316
rect 8172 28256 8236 28260
rect 8252 28316 8316 28320
rect 8252 28260 8256 28316
rect 8256 28260 8312 28316
rect 8312 28260 8316 28316
rect 8252 28256 8316 28260
rect 2352 27772 2416 27776
rect 2352 27716 2356 27772
rect 2356 27716 2412 27772
rect 2412 27716 2416 27772
rect 2352 27712 2416 27716
rect 2432 27772 2496 27776
rect 2432 27716 2436 27772
rect 2436 27716 2492 27772
rect 2492 27716 2496 27772
rect 2432 27712 2496 27716
rect 2512 27772 2576 27776
rect 2512 27716 2516 27772
rect 2516 27716 2572 27772
rect 2572 27716 2576 27772
rect 2512 27712 2576 27716
rect 2592 27772 2656 27776
rect 2592 27716 2596 27772
rect 2596 27716 2652 27772
rect 2652 27716 2656 27772
rect 2592 27712 2656 27716
rect 7352 27772 7416 27776
rect 7352 27716 7356 27772
rect 7356 27716 7412 27772
rect 7412 27716 7416 27772
rect 7352 27712 7416 27716
rect 7432 27772 7496 27776
rect 7432 27716 7436 27772
rect 7436 27716 7492 27772
rect 7492 27716 7496 27772
rect 7432 27712 7496 27716
rect 7512 27772 7576 27776
rect 7512 27716 7516 27772
rect 7516 27716 7572 27772
rect 7572 27716 7576 27772
rect 7512 27712 7576 27716
rect 7592 27772 7656 27776
rect 7592 27716 7596 27772
rect 7596 27716 7652 27772
rect 7652 27716 7656 27772
rect 7592 27712 7656 27716
rect 3012 27228 3076 27232
rect 3012 27172 3016 27228
rect 3016 27172 3072 27228
rect 3072 27172 3076 27228
rect 3012 27168 3076 27172
rect 3092 27228 3156 27232
rect 3092 27172 3096 27228
rect 3096 27172 3152 27228
rect 3152 27172 3156 27228
rect 3092 27168 3156 27172
rect 3172 27228 3236 27232
rect 3172 27172 3176 27228
rect 3176 27172 3232 27228
rect 3232 27172 3236 27228
rect 3172 27168 3236 27172
rect 3252 27228 3316 27232
rect 3252 27172 3256 27228
rect 3256 27172 3312 27228
rect 3312 27172 3316 27228
rect 3252 27168 3316 27172
rect 8012 27228 8076 27232
rect 8012 27172 8016 27228
rect 8016 27172 8072 27228
rect 8072 27172 8076 27228
rect 8012 27168 8076 27172
rect 8092 27228 8156 27232
rect 8092 27172 8096 27228
rect 8096 27172 8152 27228
rect 8152 27172 8156 27228
rect 8092 27168 8156 27172
rect 8172 27228 8236 27232
rect 8172 27172 8176 27228
rect 8176 27172 8232 27228
rect 8232 27172 8236 27228
rect 8172 27168 8236 27172
rect 8252 27228 8316 27232
rect 8252 27172 8256 27228
rect 8256 27172 8312 27228
rect 8312 27172 8316 27228
rect 8252 27168 8316 27172
rect 2352 26684 2416 26688
rect 2352 26628 2356 26684
rect 2356 26628 2412 26684
rect 2412 26628 2416 26684
rect 2352 26624 2416 26628
rect 2432 26684 2496 26688
rect 2432 26628 2436 26684
rect 2436 26628 2492 26684
rect 2492 26628 2496 26684
rect 2432 26624 2496 26628
rect 2512 26684 2576 26688
rect 2512 26628 2516 26684
rect 2516 26628 2572 26684
rect 2572 26628 2576 26684
rect 2512 26624 2576 26628
rect 2592 26684 2656 26688
rect 2592 26628 2596 26684
rect 2596 26628 2652 26684
rect 2652 26628 2656 26684
rect 2592 26624 2656 26628
rect 7352 26684 7416 26688
rect 7352 26628 7356 26684
rect 7356 26628 7412 26684
rect 7412 26628 7416 26684
rect 7352 26624 7416 26628
rect 7432 26684 7496 26688
rect 7432 26628 7436 26684
rect 7436 26628 7492 26684
rect 7492 26628 7496 26684
rect 7432 26624 7496 26628
rect 7512 26684 7576 26688
rect 7512 26628 7516 26684
rect 7516 26628 7572 26684
rect 7572 26628 7576 26684
rect 7512 26624 7576 26628
rect 7592 26684 7656 26688
rect 7592 26628 7596 26684
rect 7596 26628 7652 26684
rect 7652 26628 7656 26684
rect 7592 26624 7656 26628
rect 3012 26140 3076 26144
rect 3012 26084 3016 26140
rect 3016 26084 3072 26140
rect 3072 26084 3076 26140
rect 3012 26080 3076 26084
rect 3092 26140 3156 26144
rect 3092 26084 3096 26140
rect 3096 26084 3152 26140
rect 3152 26084 3156 26140
rect 3092 26080 3156 26084
rect 3172 26140 3236 26144
rect 3172 26084 3176 26140
rect 3176 26084 3232 26140
rect 3232 26084 3236 26140
rect 3172 26080 3236 26084
rect 3252 26140 3316 26144
rect 3252 26084 3256 26140
rect 3256 26084 3312 26140
rect 3312 26084 3316 26140
rect 3252 26080 3316 26084
rect 8012 26140 8076 26144
rect 8012 26084 8016 26140
rect 8016 26084 8072 26140
rect 8072 26084 8076 26140
rect 8012 26080 8076 26084
rect 8092 26140 8156 26144
rect 8092 26084 8096 26140
rect 8096 26084 8152 26140
rect 8152 26084 8156 26140
rect 8092 26080 8156 26084
rect 8172 26140 8236 26144
rect 8172 26084 8176 26140
rect 8176 26084 8232 26140
rect 8232 26084 8236 26140
rect 8172 26080 8236 26084
rect 8252 26140 8316 26144
rect 8252 26084 8256 26140
rect 8256 26084 8312 26140
rect 8312 26084 8316 26140
rect 8252 26080 8316 26084
rect 2352 25596 2416 25600
rect 2352 25540 2356 25596
rect 2356 25540 2412 25596
rect 2412 25540 2416 25596
rect 2352 25536 2416 25540
rect 2432 25596 2496 25600
rect 2432 25540 2436 25596
rect 2436 25540 2492 25596
rect 2492 25540 2496 25596
rect 2432 25536 2496 25540
rect 2512 25596 2576 25600
rect 2512 25540 2516 25596
rect 2516 25540 2572 25596
rect 2572 25540 2576 25596
rect 2512 25536 2576 25540
rect 2592 25596 2656 25600
rect 2592 25540 2596 25596
rect 2596 25540 2652 25596
rect 2652 25540 2656 25596
rect 2592 25536 2656 25540
rect 7352 25596 7416 25600
rect 7352 25540 7356 25596
rect 7356 25540 7412 25596
rect 7412 25540 7416 25596
rect 7352 25536 7416 25540
rect 7432 25596 7496 25600
rect 7432 25540 7436 25596
rect 7436 25540 7492 25596
rect 7492 25540 7496 25596
rect 7432 25536 7496 25540
rect 7512 25596 7576 25600
rect 7512 25540 7516 25596
rect 7516 25540 7572 25596
rect 7572 25540 7576 25596
rect 7512 25536 7576 25540
rect 7592 25596 7656 25600
rect 7592 25540 7596 25596
rect 7596 25540 7652 25596
rect 7652 25540 7656 25596
rect 7592 25536 7656 25540
rect 3012 25052 3076 25056
rect 3012 24996 3016 25052
rect 3016 24996 3072 25052
rect 3072 24996 3076 25052
rect 3012 24992 3076 24996
rect 3092 25052 3156 25056
rect 3092 24996 3096 25052
rect 3096 24996 3152 25052
rect 3152 24996 3156 25052
rect 3092 24992 3156 24996
rect 3172 25052 3236 25056
rect 3172 24996 3176 25052
rect 3176 24996 3232 25052
rect 3232 24996 3236 25052
rect 3172 24992 3236 24996
rect 3252 25052 3316 25056
rect 3252 24996 3256 25052
rect 3256 24996 3312 25052
rect 3312 24996 3316 25052
rect 3252 24992 3316 24996
rect 8012 25052 8076 25056
rect 8012 24996 8016 25052
rect 8016 24996 8072 25052
rect 8072 24996 8076 25052
rect 8012 24992 8076 24996
rect 8092 25052 8156 25056
rect 8092 24996 8096 25052
rect 8096 24996 8152 25052
rect 8152 24996 8156 25052
rect 8092 24992 8156 24996
rect 8172 25052 8236 25056
rect 8172 24996 8176 25052
rect 8176 24996 8232 25052
rect 8232 24996 8236 25052
rect 8172 24992 8236 24996
rect 8252 25052 8316 25056
rect 8252 24996 8256 25052
rect 8256 24996 8312 25052
rect 8312 24996 8316 25052
rect 8252 24992 8316 24996
rect 2352 24508 2416 24512
rect 2352 24452 2356 24508
rect 2356 24452 2412 24508
rect 2412 24452 2416 24508
rect 2352 24448 2416 24452
rect 2432 24508 2496 24512
rect 2432 24452 2436 24508
rect 2436 24452 2492 24508
rect 2492 24452 2496 24508
rect 2432 24448 2496 24452
rect 2512 24508 2576 24512
rect 2512 24452 2516 24508
rect 2516 24452 2572 24508
rect 2572 24452 2576 24508
rect 2512 24448 2576 24452
rect 2592 24508 2656 24512
rect 2592 24452 2596 24508
rect 2596 24452 2652 24508
rect 2652 24452 2656 24508
rect 2592 24448 2656 24452
rect 7352 24508 7416 24512
rect 7352 24452 7356 24508
rect 7356 24452 7412 24508
rect 7412 24452 7416 24508
rect 7352 24448 7416 24452
rect 7432 24508 7496 24512
rect 7432 24452 7436 24508
rect 7436 24452 7492 24508
rect 7492 24452 7496 24508
rect 7432 24448 7496 24452
rect 7512 24508 7576 24512
rect 7512 24452 7516 24508
rect 7516 24452 7572 24508
rect 7572 24452 7576 24508
rect 7512 24448 7576 24452
rect 7592 24508 7656 24512
rect 7592 24452 7596 24508
rect 7596 24452 7652 24508
rect 7652 24452 7656 24508
rect 7592 24448 7656 24452
rect 3012 23964 3076 23968
rect 3012 23908 3016 23964
rect 3016 23908 3072 23964
rect 3072 23908 3076 23964
rect 3012 23904 3076 23908
rect 3092 23964 3156 23968
rect 3092 23908 3096 23964
rect 3096 23908 3152 23964
rect 3152 23908 3156 23964
rect 3092 23904 3156 23908
rect 3172 23964 3236 23968
rect 3172 23908 3176 23964
rect 3176 23908 3232 23964
rect 3232 23908 3236 23964
rect 3172 23904 3236 23908
rect 3252 23964 3316 23968
rect 3252 23908 3256 23964
rect 3256 23908 3312 23964
rect 3312 23908 3316 23964
rect 3252 23904 3316 23908
rect 8012 23964 8076 23968
rect 8012 23908 8016 23964
rect 8016 23908 8072 23964
rect 8072 23908 8076 23964
rect 8012 23904 8076 23908
rect 8092 23964 8156 23968
rect 8092 23908 8096 23964
rect 8096 23908 8152 23964
rect 8152 23908 8156 23964
rect 8092 23904 8156 23908
rect 8172 23964 8236 23968
rect 8172 23908 8176 23964
rect 8176 23908 8232 23964
rect 8232 23908 8236 23964
rect 8172 23904 8236 23908
rect 8252 23964 8316 23968
rect 8252 23908 8256 23964
rect 8256 23908 8312 23964
rect 8312 23908 8316 23964
rect 8252 23904 8316 23908
rect 2352 23420 2416 23424
rect 2352 23364 2356 23420
rect 2356 23364 2412 23420
rect 2412 23364 2416 23420
rect 2352 23360 2416 23364
rect 2432 23420 2496 23424
rect 2432 23364 2436 23420
rect 2436 23364 2492 23420
rect 2492 23364 2496 23420
rect 2432 23360 2496 23364
rect 2512 23420 2576 23424
rect 2512 23364 2516 23420
rect 2516 23364 2572 23420
rect 2572 23364 2576 23420
rect 2512 23360 2576 23364
rect 2592 23420 2656 23424
rect 2592 23364 2596 23420
rect 2596 23364 2652 23420
rect 2652 23364 2656 23420
rect 2592 23360 2656 23364
rect 7352 23420 7416 23424
rect 7352 23364 7356 23420
rect 7356 23364 7412 23420
rect 7412 23364 7416 23420
rect 7352 23360 7416 23364
rect 7432 23420 7496 23424
rect 7432 23364 7436 23420
rect 7436 23364 7492 23420
rect 7492 23364 7496 23420
rect 7432 23360 7496 23364
rect 7512 23420 7576 23424
rect 7512 23364 7516 23420
rect 7516 23364 7572 23420
rect 7572 23364 7576 23420
rect 7512 23360 7576 23364
rect 7592 23420 7656 23424
rect 7592 23364 7596 23420
rect 7596 23364 7652 23420
rect 7652 23364 7656 23420
rect 7592 23360 7656 23364
rect 3012 22876 3076 22880
rect 3012 22820 3016 22876
rect 3016 22820 3072 22876
rect 3072 22820 3076 22876
rect 3012 22816 3076 22820
rect 3092 22876 3156 22880
rect 3092 22820 3096 22876
rect 3096 22820 3152 22876
rect 3152 22820 3156 22876
rect 3092 22816 3156 22820
rect 3172 22876 3236 22880
rect 3172 22820 3176 22876
rect 3176 22820 3232 22876
rect 3232 22820 3236 22876
rect 3172 22816 3236 22820
rect 3252 22876 3316 22880
rect 3252 22820 3256 22876
rect 3256 22820 3312 22876
rect 3312 22820 3316 22876
rect 3252 22816 3316 22820
rect 8012 22876 8076 22880
rect 8012 22820 8016 22876
rect 8016 22820 8072 22876
rect 8072 22820 8076 22876
rect 8012 22816 8076 22820
rect 8092 22876 8156 22880
rect 8092 22820 8096 22876
rect 8096 22820 8152 22876
rect 8152 22820 8156 22876
rect 8092 22816 8156 22820
rect 8172 22876 8236 22880
rect 8172 22820 8176 22876
rect 8176 22820 8232 22876
rect 8232 22820 8236 22876
rect 8172 22816 8236 22820
rect 8252 22876 8316 22880
rect 8252 22820 8256 22876
rect 8256 22820 8312 22876
rect 8312 22820 8316 22876
rect 8252 22816 8316 22820
rect 2352 22332 2416 22336
rect 2352 22276 2356 22332
rect 2356 22276 2412 22332
rect 2412 22276 2416 22332
rect 2352 22272 2416 22276
rect 2432 22332 2496 22336
rect 2432 22276 2436 22332
rect 2436 22276 2492 22332
rect 2492 22276 2496 22332
rect 2432 22272 2496 22276
rect 2512 22332 2576 22336
rect 2512 22276 2516 22332
rect 2516 22276 2572 22332
rect 2572 22276 2576 22332
rect 2512 22272 2576 22276
rect 2592 22332 2656 22336
rect 2592 22276 2596 22332
rect 2596 22276 2652 22332
rect 2652 22276 2656 22332
rect 2592 22272 2656 22276
rect 7352 22332 7416 22336
rect 7352 22276 7356 22332
rect 7356 22276 7412 22332
rect 7412 22276 7416 22332
rect 7352 22272 7416 22276
rect 7432 22332 7496 22336
rect 7432 22276 7436 22332
rect 7436 22276 7492 22332
rect 7492 22276 7496 22332
rect 7432 22272 7496 22276
rect 7512 22332 7576 22336
rect 7512 22276 7516 22332
rect 7516 22276 7572 22332
rect 7572 22276 7576 22332
rect 7512 22272 7576 22276
rect 7592 22332 7656 22336
rect 7592 22276 7596 22332
rect 7596 22276 7652 22332
rect 7652 22276 7656 22332
rect 7592 22272 7656 22276
rect 3012 21788 3076 21792
rect 3012 21732 3016 21788
rect 3016 21732 3072 21788
rect 3072 21732 3076 21788
rect 3012 21728 3076 21732
rect 3092 21788 3156 21792
rect 3092 21732 3096 21788
rect 3096 21732 3152 21788
rect 3152 21732 3156 21788
rect 3092 21728 3156 21732
rect 3172 21788 3236 21792
rect 3172 21732 3176 21788
rect 3176 21732 3232 21788
rect 3232 21732 3236 21788
rect 3172 21728 3236 21732
rect 3252 21788 3316 21792
rect 3252 21732 3256 21788
rect 3256 21732 3312 21788
rect 3312 21732 3316 21788
rect 3252 21728 3316 21732
rect 8012 21788 8076 21792
rect 8012 21732 8016 21788
rect 8016 21732 8072 21788
rect 8072 21732 8076 21788
rect 8012 21728 8076 21732
rect 8092 21788 8156 21792
rect 8092 21732 8096 21788
rect 8096 21732 8152 21788
rect 8152 21732 8156 21788
rect 8092 21728 8156 21732
rect 8172 21788 8236 21792
rect 8172 21732 8176 21788
rect 8176 21732 8232 21788
rect 8232 21732 8236 21788
rect 8172 21728 8236 21732
rect 8252 21788 8316 21792
rect 8252 21732 8256 21788
rect 8256 21732 8312 21788
rect 8312 21732 8316 21788
rect 8252 21728 8316 21732
rect 2352 21244 2416 21248
rect 2352 21188 2356 21244
rect 2356 21188 2412 21244
rect 2412 21188 2416 21244
rect 2352 21184 2416 21188
rect 2432 21244 2496 21248
rect 2432 21188 2436 21244
rect 2436 21188 2492 21244
rect 2492 21188 2496 21244
rect 2432 21184 2496 21188
rect 2512 21244 2576 21248
rect 2512 21188 2516 21244
rect 2516 21188 2572 21244
rect 2572 21188 2576 21244
rect 2512 21184 2576 21188
rect 2592 21244 2656 21248
rect 2592 21188 2596 21244
rect 2596 21188 2652 21244
rect 2652 21188 2656 21244
rect 2592 21184 2656 21188
rect 7352 21244 7416 21248
rect 7352 21188 7356 21244
rect 7356 21188 7412 21244
rect 7412 21188 7416 21244
rect 7352 21184 7416 21188
rect 7432 21244 7496 21248
rect 7432 21188 7436 21244
rect 7436 21188 7492 21244
rect 7492 21188 7496 21244
rect 7432 21184 7496 21188
rect 7512 21244 7576 21248
rect 7512 21188 7516 21244
rect 7516 21188 7572 21244
rect 7572 21188 7576 21244
rect 7512 21184 7576 21188
rect 7592 21244 7656 21248
rect 7592 21188 7596 21244
rect 7596 21188 7652 21244
rect 7652 21188 7656 21244
rect 7592 21184 7656 21188
rect 3012 20700 3076 20704
rect 3012 20644 3016 20700
rect 3016 20644 3072 20700
rect 3072 20644 3076 20700
rect 3012 20640 3076 20644
rect 3092 20700 3156 20704
rect 3092 20644 3096 20700
rect 3096 20644 3152 20700
rect 3152 20644 3156 20700
rect 3092 20640 3156 20644
rect 3172 20700 3236 20704
rect 3172 20644 3176 20700
rect 3176 20644 3232 20700
rect 3232 20644 3236 20700
rect 3172 20640 3236 20644
rect 3252 20700 3316 20704
rect 3252 20644 3256 20700
rect 3256 20644 3312 20700
rect 3312 20644 3316 20700
rect 3252 20640 3316 20644
rect 8012 20700 8076 20704
rect 8012 20644 8016 20700
rect 8016 20644 8072 20700
rect 8072 20644 8076 20700
rect 8012 20640 8076 20644
rect 8092 20700 8156 20704
rect 8092 20644 8096 20700
rect 8096 20644 8152 20700
rect 8152 20644 8156 20700
rect 8092 20640 8156 20644
rect 8172 20700 8236 20704
rect 8172 20644 8176 20700
rect 8176 20644 8232 20700
rect 8232 20644 8236 20700
rect 8172 20640 8236 20644
rect 8252 20700 8316 20704
rect 8252 20644 8256 20700
rect 8256 20644 8312 20700
rect 8312 20644 8316 20700
rect 8252 20640 8316 20644
rect 2352 20156 2416 20160
rect 2352 20100 2356 20156
rect 2356 20100 2412 20156
rect 2412 20100 2416 20156
rect 2352 20096 2416 20100
rect 2432 20156 2496 20160
rect 2432 20100 2436 20156
rect 2436 20100 2492 20156
rect 2492 20100 2496 20156
rect 2432 20096 2496 20100
rect 2512 20156 2576 20160
rect 2512 20100 2516 20156
rect 2516 20100 2572 20156
rect 2572 20100 2576 20156
rect 2512 20096 2576 20100
rect 2592 20156 2656 20160
rect 2592 20100 2596 20156
rect 2596 20100 2652 20156
rect 2652 20100 2656 20156
rect 2592 20096 2656 20100
rect 7352 20156 7416 20160
rect 7352 20100 7356 20156
rect 7356 20100 7412 20156
rect 7412 20100 7416 20156
rect 7352 20096 7416 20100
rect 7432 20156 7496 20160
rect 7432 20100 7436 20156
rect 7436 20100 7492 20156
rect 7492 20100 7496 20156
rect 7432 20096 7496 20100
rect 7512 20156 7576 20160
rect 7512 20100 7516 20156
rect 7516 20100 7572 20156
rect 7572 20100 7576 20156
rect 7512 20096 7576 20100
rect 7592 20156 7656 20160
rect 7592 20100 7596 20156
rect 7596 20100 7652 20156
rect 7652 20100 7656 20156
rect 7592 20096 7656 20100
rect 3012 19612 3076 19616
rect 3012 19556 3016 19612
rect 3016 19556 3072 19612
rect 3072 19556 3076 19612
rect 3012 19552 3076 19556
rect 3092 19612 3156 19616
rect 3092 19556 3096 19612
rect 3096 19556 3152 19612
rect 3152 19556 3156 19612
rect 3092 19552 3156 19556
rect 3172 19612 3236 19616
rect 3172 19556 3176 19612
rect 3176 19556 3232 19612
rect 3232 19556 3236 19612
rect 3172 19552 3236 19556
rect 3252 19612 3316 19616
rect 3252 19556 3256 19612
rect 3256 19556 3312 19612
rect 3312 19556 3316 19612
rect 3252 19552 3316 19556
rect 8012 19612 8076 19616
rect 8012 19556 8016 19612
rect 8016 19556 8072 19612
rect 8072 19556 8076 19612
rect 8012 19552 8076 19556
rect 8092 19612 8156 19616
rect 8092 19556 8096 19612
rect 8096 19556 8152 19612
rect 8152 19556 8156 19612
rect 8092 19552 8156 19556
rect 8172 19612 8236 19616
rect 8172 19556 8176 19612
rect 8176 19556 8232 19612
rect 8232 19556 8236 19612
rect 8172 19552 8236 19556
rect 8252 19612 8316 19616
rect 8252 19556 8256 19612
rect 8256 19556 8312 19612
rect 8312 19556 8316 19612
rect 8252 19552 8316 19556
rect 2352 19068 2416 19072
rect 2352 19012 2356 19068
rect 2356 19012 2412 19068
rect 2412 19012 2416 19068
rect 2352 19008 2416 19012
rect 2432 19068 2496 19072
rect 2432 19012 2436 19068
rect 2436 19012 2492 19068
rect 2492 19012 2496 19068
rect 2432 19008 2496 19012
rect 2512 19068 2576 19072
rect 2512 19012 2516 19068
rect 2516 19012 2572 19068
rect 2572 19012 2576 19068
rect 2512 19008 2576 19012
rect 2592 19068 2656 19072
rect 2592 19012 2596 19068
rect 2596 19012 2652 19068
rect 2652 19012 2656 19068
rect 2592 19008 2656 19012
rect 7352 19068 7416 19072
rect 7352 19012 7356 19068
rect 7356 19012 7412 19068
rect 7412 19012 7416 19068
rect 7352 19008 7416 19012
rect 7432 19068 7496 19072
rect 7432 19012 7436 19068
rect 7436 19012 7492 19068
rect 7492 19012 7496 19068
rect 7432 19008 7496 19012
rect 7512 19068 7576 19072
rect 7512 19012 7516 19068
rect 7516 19012 7572 19068
rect 7572 19012 7576 19068
rect 7512 19008 7576 19012
rect 7592 19068 7656 19072
rect 7592 19012 7596 19068
rect 7596 19012 7652 19068
rect 7652 19012 7656 19068
rect 7592 19008 7656 19012
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 3172 18524 3236 18528
rect 3172 18468 3176 18524
rect 3176 18468 3232 18524
rect 3232 18468 3236 18524
rect 3172 18464 3236 18468
rect 3252 18524 3316 18528
rect 3252 18468 3256 18524
rect 3256 18468 3312 18524
rect 3312 18468 3316 18524
rect 3252 18464 3316 18468
rect 8012 18524 8076 18528
rect 8012 18468 8016 18524
rect 8016 18468 8072 18524
rect 8072 18468 8076 18524
rect 8012 18464 8076 18468
rect 8092 18524 8156 18528
rect 8092 18468 8096 18524
rect 8096 18468 8152 18524
rect 8152 18468 8156 18524
rect 8092 18464 8156 18468
rect 8172 18524 8236 18528
rect 8172 18468 8176 18524
rect 8176 18468 8232 18524
rect 8232 18468 8236 18524
rect 8172 18464 8236 18468
rect 8252 18524 8316 18528
rect 8252 18468 8256 18524
rect 8256 18468 8312 18524
rect 8312 18468 8316 18524
rect 8252 18464 8316 18468
rect 2352 17980 2416 17984
rect 2352 17924 2356 17980
rect 2356 17924 2412 17980
rect 2412 17924 2416 17980
rect 2352 17920 2416 17924
rect 2432 17980 2496 17984
rect 2432 17924 2436 17980
rect 2436 17924 2492 17980
rect 2492 17924 2496 17980
rect 2432 17920 2496 17924
rect 2512 17980 2576 17984
rect 2512 17924 2516 17980
rect 2516 17924 2572 17980
rect 2572 17924 2576 17980
rect 2512 17920 2576 17924
rect 2592 17980 2656 17984
rect 2592 17924 2596 17980
rect 2596 17924 2652 17980
rect 2652 17924 2656 17980
rect 2592 17920 2656 17924
rect 7352 17980 7416 17984
rect 7352 17924 7356 17980
rect 7356 17924 7412 17980
rect 7412 17924 7416 17980
rect 7352 17920 7416 17924
rect 7432 17980 7496 17984
rect 7432 17924 7436 17980
rect 7436 17924 7492 17980
rect 7492 17924 7496 17980
rect 7432 17920 7496 17924
rect 7512 17980 7576 17984
rect 7512 17924 7516 17980
rect 7516 17924 7572 17980
rect 7572 17924 7576 17980
rect 7512 17920 7576 17924
rect 7592 17980 7656 17984
rect 7592 17924 7596 17980
rect 7596 17924 7652 17980
rect 7652 17924 7656 17980
rect 7592 17920 7656 17924
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 3172 17436 3236 17440
rect 3172 17380 3176 17436
rect 3176 17380 3232 17436
rect 3232 17380 3236 17436
rect 3172 17376 3236 17380
rect 3252 17436 3316 17440
rect 3252 17380 3256 17436
rect 3256 17380 3312 17436
rect 3312 17380 3316 17436
rect 3252 17376 3316 17380
rect 8012 17436 8076 17440
rect 8012 17380 8016 17436
rect 8016 17380 8072 17436
rect 8072 17380 8076 17436
rect 8012 17376 8076 17380
rect 8092 17436 8156 17440
rect 8092 17380 8096 17436
rect 8096 17380 8152 17436
rect 8152 17380 8156 17436
rect 8092 17376 8156 17380
rect 8172 17436 8236 17440
rect 8172 17380 8176 17436
rect 8176 17380 8232 17436
rect 8232 17380 8236 17436
rect 8172 17376 8236 17380
rect 8252 17436 8316 17440
rect 8252 17380 8256 17436
rect 8256 17380 8312 17436
rect 8312 17380 8316 17436
rect 8252 17376 8316 17380
rect 2352 16892 2416 16896
rect 2352 16836 2356 16892
rect 2356 16836 2412 16892
rect 2412 16836 2416 16892
rect 2352 16832 2416 16836
rect 2432 16892 2496 16896
rect 2432 16836 2436 16892
rect 2436 16836 2492 16892
rect 2492 16836 2496 16892
rect 2432 16832 2496 16836
rect 2512 16892 2576 16896
rect 2512 16836 2516 16892
rect 2516 16836 2572 16892
rect 2572 16836 2576 16892
rect 2512 16832 2576 16836
rect 2592 16892 2656 16896
rect 2592 16836 2596 16892
rect 2596 16836 2652 16892
rect 2652 16836 2656 16892
rect 2592 16832 2656 16836
rect 7352 16892 7416 16896
rect 7352 16836 7356 16892
rect 7356 16836 7412 16892
rect 7412 16836 7416 16892
rect 7352 16832 7416 16836
rect 7432 16892 7496 16896
rect 7432 16836 7436 16892
rect 7436 16836 7492 16892
rect 7492 16836 7496 16892
rect 7432 16832 7496 16836
rect 7512 16892 7576 16896
rect 7512 16836 7516 16892
rect 7516 16836 7572 16892
rect 7572 16836 7576 16892
rect 7512 16832 7576 16836
rect 7592 16892 7656 16896
rect 7592 16836 7596 16892
rect 7596 16836 7652 16892
rect 7652 16836 7656 16892
rect 7592 16832 7656 16836
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 3172 16348 3236 16352
rect 3172 16292 3176 16348
rect 3176 16292 3232 16348
rect 3232 16292 3236 16348
rect 3172 16288 3236 16292
rect 3252 16348 3316 16352
rect 3252 16292 3256 16348
rect 3256 16292 3312 16348
rect 3312 16292 3316 16348
rect 3252 16288 3316 16292
rect 8012 16348 8076 16352
rect 8012 16292 8016 16348
rect 8016 16292 8072 16348
rect 8072 16292 8076 16348
rect 8012 16288 8076 16292
rect 8092 16348 8156 16352
rect 8092 16292 8096 16348
rect 8096 16292 8152 16348
rect 8152 16292 8156 16348
rect 8092 16288 8156 16292
rect 8172 16348 8236 16352
rect 8172 16292 8176 16348
rect 8176 16292 8232 16348
rect 8232 16292 8236 16348
rect 8172 16288 8236 16292
rect 8252 16348 8316 16352
rect 8252 16292 8256 16348
rect 8256 16292 8312 16348
rect 8312 16292 8316 16348
rect 8252 16288 8316 16292
rect 2352 15804 2416 15808
rect 2352 15748 2356 15804
rect 2356 15748 2412 15804
rect 2412 15748 2416 15804
rect 2352 15744 2416 15748
rect 2432 15804 2496 15808
rect 2432 15748 2436 15804
rect 2436 15748 2492 15804
rect 2492 15748 2496 15804
rect 2432 15744 2496 15748
rect 2512 15804 2576 15808
rect 2512 15748 2516 15804
rect 2516 15748 2572 15804
rect 2572 15748 2576 15804
rect 2512 15744 2576 15748
rect 2592 15804 2656 15808
rect 2592 15748 2596 15804
rect 2596 15748 2652 15804
rect 2652 15748 2656 15804
rect 2592 15744 2656 15748
rect 7352 15804 7416 15808
rect 7352 15748 7356 15804
rect 7356 15748 7412 15804
rect 7412 15748 7416 15804
rect 7352 15744 7416 15748
rect 7432 15804 7496 15808
rect 7432 15748 7436 15804
rect 7436 15748 7492 15804
rect 7492 15748 7496 15804
rect 7432 15744 7496 15748
rect 7512 15804 7576 15808
rect 7512 15748 7516 15804
rect 7516 15748 7572 15804
rect 7572 15748 7576 15804
rect 7512 15744 7576 15748
rect 7592 15804 7656 15808
rect 7592 15748 7596 15804
rect 7596 15748 7652 15804
rect 7652 15748 7656 15804
rect 7592 15744 7656 15748
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 3172 15260 3236 15264
rect 3172 15204 3176 15260
rect 3176 15204 3232 15260
rect 3232 15204 3236 15260
rect 3172 15200 3236 15204
rect 3252 15260 3316 15264
rect 3252 15204 3256 15260
rect 3256 15204 3312 15260
rect 3312 15204 3316 15260
rect 3252 15200 3316 15204
rect 8012 15260 8076 15264
rect 8012 15204 8016 15260
rect 8016 15204 8072 15260
rect 8072 15204 8076 15260
rect 8012 15200 8076 15204
rect 8092 15260 8156 15264
rect 8092 15204 8096 15260
rect 8096 15204 8152 15260
rect 8152 15204 8156 15260
rect 8092 15200 8156 15204
rect 8172 15260 8236 15264
rect 8172 15204 8176 15260
rect 8176 15204 8232 15260
rect 8232 15204 8236 15260
rect 8172 15200 8236 15204
rect 8252 15260 8316 15264
rect 8252 15204 8256 15260
rect 8256 15204 8312 15260
rect 8312 15204 8316 15260
rect 8252 15200 8316 15204
rect 2352 14716 2416 14720
rect 2352 14660 2356 14716
rect 2356 14660 2412 14716
rect 2412 14660 2416 14716
rect 2352 14656 2416 14660
rect 2432 14716 2496 14720
rect 2432 14660 2436 14716
rect 2436 14660 2492 14716
rect 2492 14660 2496 14716
rect 2432 14656 2496 14660
rect 2512 14716 2576 14720
rect 2512 14660 2516 14716
rect 2516 14660 2572 14716
rect 2572 14660 2576 14716
rect 2512 14656 2576 14660
rect 2592 14716 2656 14720
rect 2592 14660 2596 14716
rect 2596 14660 2652 14716
rect 2652 14660 2656 14716
rect 2592 14656 2656 14660
rect 7352 14716 7416 14720
rect 7352 14660 7356 14716
rect 7356 14660 7412 14716
rect 7412 14660 7416 14716
rect 7352 14656 7416 14660
rect 7432 14716 7496 14720
rect 7432 14660 7436 14716
rect 7436 14660 7492 14716
rect 7492 14660 7496 14716
rect 7432 14656 7496 14660
rect 7512 14716 7576 14720
rect 7512 14660 7516 14716
rect 7516 14660 7572 14716
rect 7572 14660 7576 14716
rect 7512 14656 7576 14660
rect 7592 14716 7656 14720
rect 7592 14660 7596 14716
rect 7596 14660 7652 14716
rect 7652 14660 7656 14716
rect 7592 14656 7656 14660
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 3172 14172 3236 14176
rect 3172 14116 3176 14172
rect 3176 14116 3232 14172
rect 3232 14116 3236 14172
rect 3172 14112 3236 14116
rect 3252 14172 3316 14176
rect 3252 14116 3256 14172
rect 3256 14116 3312 14172
rect 3312 14116 3316 14172
rect 3252 14112 3316 14116
rect 8012 14172 8076 14176
rect 8012 14116 8016 14172
rect 8016 14116 8072 14172
rect 8072 14116 8076 14172
rect 8012 14112 8076 14116
rect 8092 14172 8156 14176
rect 8092 14116 8096 14172
rect 8096 14116 8152 14172
rect 8152 14116 8156 14172
rect 8092 14112 8156 14116
rect 8172 14172 8236 14176
rect 8172 14116 8176 14172
rect 8176 14116 8232 14172
rect 8232 14116 8236 14172
rect 8172 14112 8236 14116
rect 8252 14172 8316 14176
rect 8252 14116 8256 14172
rect 8256 14116 8312 14172
rect 8312 14116 8316 14172
rect 8252 14112 8316 14116
rect 2352 13628 2416 13632
rect 2352 13572 2356 13628
rect 2356 13572 2412 13628
rect 2412 13572 2416 13628
rect 2352 13568 2416 13572
rect 2432 13628 2496 13632
rect 2432 13572 2436 13628
rect 2436 13572 2492 13628
rect 2492 13572 2496 13628
rect 2432 13568 2496 13572
rect 2512 13628 2576 13632
rect 2512 13572 2516 13628
rect 2516 13572 2572 13628
rect 2572 13572 2576 13628
rect 2512 13568 2576 13572
rect 2592 13628 2656 13632
rect 2592 13572 2596 13628
rect 2596 13572 2652 13628
rect 2652 13572 2656 13628
rect 2592 13568 2656 13572
rect 7352 13628 7416 13632
rect 7352 13572 7356 13628
rect 7356 13572 7412 13628
rect 7412 13572 7416 13628
rect 7352 13568 7416 13572
rect 7432 13628 7496 13632
rect 7432 13572 7436 13628
rect 7436 13572 7492 13628
rect 7492 13572 7496 13628
rect 7432 13568 7496 13572
rect 7512 13628 7576 13632
rect 7512 13572 7516 13628
rect 7516 13572 7572 13628
rect 7572 13572 7576 13628
rect 7512 13568 7576 13572
rect 7592 13628 7656 13632
rect 7592 13572 7596 13628
rect 7596 13572 7652 13628
rect 7652 13572 7656 13628
rect 7592 13568 7656 13572
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 3172 13084 3236 13088
rect 3172 13028 3176 13084
rect 3176 13028 3232 13084
rect 3232 13028 3236 13084
rect 3172 13024 3236 13028
rect 3252 13084 3316 13088
rect 3252 13028 3256 13084
rect 3256 13028 3312 13084
rect 3312 13028 3316 13084
rect 3252 13024 3316 13028
rect 8012 13084 8076 13088
rect 8012 13028 8016 13084
rect 8016 13028 8072 13084
rect 8072 13028 8076 13084
rect 8012 13024 8076 13028
rect 8092 13084 8156 13088
rect 8092 13028 8096 13084
rect 8096 13028 8152 13084
rect 8152 13028 8156 13084
rect 8092 13024 8156 13028
rect 8172 13084 8236 13088
rect 8172 13028 8176 13084
rect 8176 13028 8232 13084
rect 8232 13028 8236 13084
rect 8172 13024 8236 13028
rect 8252 13084 8316 13088
rect 8252 13028 8256 13084
rect 8256 13028 8312 13084
rect 8312 13028 8316 13084
rect 8252 13024 8316 13028
rect 2352 12540 2416 12544
rect 2352 12484 2356 12540
rect 2356 12484 2412 12540
rect 2412 12484 2416 12540
rect 2352 12480 2416 12484
rect 2432 12540 2496 12544
rect 2432 12484 2436 12540
rect 2436 12484 2492 12540
rect 2492 12484 2496 12540
rect 2432 12480 2496 12484
rect 2512 12540 2576 12544
rect 2512 12484 2516 12540
rect 2516 12484 2572 12540
rect 2572 12484 2576 12540
rect 2512 12480 2576 12484
rect 2592 12540 2656 12544
rect 2592 12484 2596 12540
rect 2596 12484 2652 12540
rect 2652 12484 2656 12540
rect 2592 12480 2656 12484
rect 7352 12540 7416 12544
rect 7352 12484 7356 12540
rect 7356 12484 7412 12540
rect 7412 12484 7416 12540
rect 7352 12480 7416 12484
rect 7432 12540 7496 12544
rect 7432 12484 7436 12540
rect 7436 12484 7492 12540
rect 7492 12484 7496 12540
rect 7432 12480 7496 12484
rect 7512 12540 7576 12544
rect 7512 12484 7516 12540
rect 7516 12484 7572 12540
rect 7572 12484 7576 12540
rect 7512 12480 7576 12484
rect 7592 12540 7656 12544
rect 7592 12484 7596 12540
rect 7596 12484 7652 12540
rect 7652 12484 7656 12540
rect 7592 12480 7656 12484
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 3172 11996 3236 12000
rect 3172 11940 3176 11996
rect 3176 11940 3232 11996
rect 3232 11940 3236 11996
rect 3172 11936 3236 11940
rect 3252 11996 3316 12000
rect 3252 11940 3256 11996
rect 3256 11940 3312 11996
rect 3312 11940 3316 11996
rect 3252 11936 3316 11940
rect 8012 11996 8076 12000
rect 8012 11940 8016 11996
rect 8016 11940 8072 11996
rect 8072 11940 8076 11996
rect 8012 11936 8076 11940
rect 8092 11996 8156 12000
rect 8092 11940 8096 11996
rect 8096 11940 8152 11996
rect 8152 11940 8156 11996
rect 8092 11936 8156 11940
rect 8172 11996 8236 12000
rect 8172 11940 8176 11996
rect 8176 11940 8232 11996
rect 8232 11940 8236 11996
rect 8172 11936 8236 11940
rect 8252 11996 8316 12000
rect 8252 11940 8256 11996
rect 8256 11940 8312 11996
rect 8312 11940 8316 11996
rect 8252 11936 8316 11940
rect 2352 11452 2416 11456
rect 2352 11396 2356 11452
rect 2356 11396 2412 11452
rect 2412 11396 2416 11452
rect 2352 11392 2416 11396
rect 2432 11452 2496 11456
rect 2432 11396 2436 11452
rect 2436 11396 2492 11452
rect 2492 11396 2496 11452
rect 2432 11392 2496 11396
rect 2512 11452 2576 11456
rect 2512 11396 2516 11452
rect 2516 11396 2572 11452
rect 2572 11396 2576 11452
rect 2512 11392 2576 11396
rect 2592 11452 2656 11456
rect 2592 11396 2596 11452
rect 2596 11396 2652 11452
rect 2652 11396 2656 11452
rect 2592 11392 2656 11396
rect 7352 11452 7416 11456
rect 7352 11396 7356 11452
rect 7356 11396 7412 11452
rect 7412 11396 7416 11452
rect 7352 11392 7416 11396
rect 7432 11452 7496 11456
rect 7432 11396 7436 11452
rect 7436 11396 7492 11452
rect 7492 11396 7496 11452
rect 7432 11392 7496 11396
rect 7512 11452 7576 11456
rect 7512 11396 7516 11452
rect 7516 11396 7572 11452
rect 7572 11396 7576 11452
rect 7512 11392 7576 11396
rect 7592 11452 7656 11456
rect 7592 11396 7596 11452
rect 7596 11396 7652 11452
rect 7652 11396 7656 11452
rect 7592 11392 7656 11396
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 3172 10908 3236 10912
rect 3172 10852 3176 10908
rect 3176 10852 3232 10908
rect 3232 10852 3236 10908
rect 3172 10848 3236 10852
rect 3252 10908 3316 10912
rect 3252 10852 3256 10908
rect 3256 10852 3312 10908
rect 3312 10852 3316 10908
rect 3252 10848 3316 10852
rect 8012 10908 8076 10912
rect 8012 10852 8016 10908
rect 8016 10852 8072 10908
rect 8072 10852 8076 10908
rect 8012 10848 8076 10852
rect 8092 10908 8156 10912
rect 8092 10852 8096 10908
rect 8096 10852 8152 10908
rect 8152 10852 8156 10908
rect 8092 10848 8156 10852
rect 8172 10908 8236 10912
rect 8172 10852 8176 10908
rect 8176 10852 8232 10908
rect 8232 10852 8236 10908
rect 8172 10848 8236 10852
rect 8252 10908 8316 10912
rect 8252 10852 8256 10908
rect 8256 10852 8312 10908
rect 8312 10852 8316 10908
rect 8252 10848 8316 10852
rect 2352 10364 2416 10368
rect 2352 10308 2356 10364
rect 2356 10308 2412 10364
rect 2412 10308 2416 10364
rect 2352 10304 2416 10308
rect 2432 10364 2496 10368
rect 2432 10308 2436 10364
rect 2436 10308 2492 10364
rect 2492 10308 2496 10364
rect 2432 10304 2496 10308
rect 2512 10364 2576 10368
rect 2512 10308 2516 10364
rect 2516 10308 2572 10364
rect 2572 10308 2576 10364
rect 2512 10304 2576 10308
rect 2592 10364 2656 10368
rect 2592 10308 2596 10364
rect 2596 10308 2652 10364
rect 2652 10308 2656 10364
rect 2592 10304 2656 10308
rect 7352 10364 7416 10368
rect 7352 10308 7356 10364
rect 7356 10308 7412 10364
rect 7412 10308 7416 10364
rect 7352 10304 7416 10308
rect 7432 10364 7496 10368
rect 7432 10308 7436 10364
rect 7436 10308 7492 10364
rect 7492 10308 7496 10364
rect 7432 10304 7496 10308
rect 7512 10364 7576 10368
rect 7512 10308 7516 10364
rect 7516 10308 7572 10364
rect 7572 10308 7576 10364
rect 7512 10304 7576 10308
rect 7592 10364 7656 10368
rect 7592 10308 7596 10364
rect 7596 10308 7652 10364
rect 7652 10308 7656 10364
rect 7592 10304 7656 10308
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 3172 9820 3236 9824
rect 3172 9764 3176 9820
rect 3176 9764 3232 9820
rect 3232 9764 3236 9820
rect 3172 9760 3236 9764
rect 3252 9820 3316 9824
rect 3252 9764 3256 9820
rect 3256 9764 3312 9820
rect 3312 9764 3316 9820
rect 3252 9760 3316 9764
rect 8012 9820 8076 9824
rect 8012 9764 8016 9820
rect 8016 9764 8072 9820
rect 8072 9764 8076 9820
rect 8012 9760 8076 9764
rect 8092 9820 8156 9824
rect 8092 9764 8096 9820
rect 8096 9764 8152 9820
rect 8152 9764 8156 9820
rect 8092 9760 8156 9764
rect 8172 9820 8236 9824
rect 8172 9764 8176 9820
rect 8176 9764 8232 9820
rect 8232 9764 8236 9820
rect 8172 9760 8236 9764
rect 8252 9820 8316 9824
rect 8252 9764 8256 9820
rect 8256 9764 8312 9820
rect 8312 9764 8316 9820
rect 8252 9760 8316 9764
rect 2352 9276 2416 9280
rect 2352 9220 2356 9276
rect 2356 9220 2412 9276
rect 2412 9220 2416 9276
rect 2352 9216 2416 9220
rect 2432 9276 2496 9280
rect 2432 9220 2436 9276
rect 2436 9220 2492 9276
rect 2492 9220 2496 9276
rect 2432 9216 2496 9220
rect 2512 9276 2576 9280
rect 2512 9220 2516 9276
rect 2516 9220 2572 9276
rect 2572 9220 2576 9276
rect 2512 9216 2576 9220
rect 2592 9276 2656 9280
rect 2592 9220 2596 9276
rect 2596 9220 2652 9276
rect 2652 9220 2656 9276
rect 2592 9216 2656 9220
rect 7352 9276 7416 9280
rect 7352 9220 7356 9276
rect 7356 9220 7412 9276
rect 7412 9220 7416 9276
rect 7352 9216 7416 9220
rect 7432 9276 7496 9280
rect 7432 9220 7436 9276
rect 7436 9220 7492 9276
rect 7492 9220 7496 9276
rect 7432 9216 7496 9220
rect 7512 9276 7576 9280
rect 7512 9220 7516 9276
rect 7516 9220 7572 9276
rect 7572 9220 7576 9276
rect 7512 9216 7576 9220
rect 7592 9276 7656 9280
rect 7592 9220 7596 9276
rect 7596 9220 7652 9276
rect 7652 9220 7656 9276
rect 7592 9216 7656 9220
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 8012 8732 8076 8736
rect 8012 8676 8016 8732
rect 8016 8676 8072 8732
rect 8072 8676 8076 8732
rect 8012 8672 8076 8676
rect 8092 8732 8156 8736
rect 8092 8676 8096 8732
rect 8096 8676 8152 8732
rect 8152 8676 8156 8732
rect 8092 8672 8156 8676
rect 8172 8732 8236 8736
rect 8172 8676 8176 8732
rect 8176 8676 8232 8732
rect 8232 8676 8236 8732
rect 8172 8672 8236 8676
rect 8252 8732 8316 8736
rect 8252 8676 8256 8732
rect 8256 8676 8312 8732
rect 8312 8676 8316 8732
rect 8252 8672 8316 8676
rect 2352 8188 2416 8192
rect 2352 8132 2356 8188
rect 2356 8132 2412 8188
rect 2412 8132 2416 8188
rect 2352 8128 2416 8132
rect 2432 8188 2496 8192
rect 2432 8132 2436 8188
rect 2436 8132 2492 8188
rect 2492 8132 2496 8188
rect 2432 8128 2496 8132
rect 2512 8188 2576 8192
rect 2512 8132 2516 8188
rect 2516 8132 2572 8188
rect 2572 8132 2576 8188
rect 2512 8128 2576 8132
rect 2592 8188 2656 8192
rect 2592 8132 2596 8188
rect 2596 8132 2652 8188
rect 2652 8132 2656 8188
rect 2592 8128 2656 8132
rect 7352 8188 7416 8192
rect 7352 8132 7356 8188
rect 7356 8132 7412 8188
rect 7412 8132 7416 8188
rect 7352 8128 7416 8132
rect 7432 8188 7496 8192
rect 7432 8132 7436 8188
rect 7436 8132 7492 8188
rect 7492 8132 7496 8188
rect 7432 8128 7496 8132
rect 7512 8188 7576 8192
rect 7512 8132 7516 8188
rect 7516 8132 7572 8188
rect 7572 8132 7576 8188
rect 7512 8128 7576 8132
rect 7592 8188 7656 8192
rect 7592 8132 7596 8188
rect 7596 8132 7652 8188
rect 7652 8132 7656 8188
rect 7592 8128 7656 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 8012 7644 8076 7648
rect 8012 7588 8016 7644
rect 8016 7588 8072 7644
rect 8072 7588 8076 7644
rect 8012 7584 8076 7588
rect 8092 7644 8156 7648
rect 8092 7588 8096 7644
rect 8096 7588 8152 7644
rect 8152 7588 8156 7644
rect 8092 7584 8156 7588
rect 8172 7644 8236 7648
rect 8172 7588 8176 7644
rect 8176 7588 8232 7644
rect 8232 7588 8236 7644
rect 8172 7584 8236 7588
rect 8252 7644 8316 7648
rect 8252 7588 8256 7644
rect 8256 7588 8312 7644
rect 8312 7588 8316 7644
rect 8252 7584 8316 7588
rect 2352 7100 2416 7104
rect 2352 7044 2356 7100
rect 2356 7044 2412 7100
rect 2412 7044 2416 7100
rect 2352 7040 2416 7044
rect 2432 7100 2496 7104
rect 2432 7044 2436 7100
rect 2436 7044 2492 7100
rect 2492 7044 2496 7100
rect 2432 7040 2496 7044
rect 2512 7100 2576 7104
rect 2512 7044 2516 7100
rect 2516 7044 2572 7100
rect 2572 7044 2576 7100
rect 2512 7040 2576 7044
rect 2592 7100 2656 7104
rect 2592 7044 2596 7100
rect 2596 7044 2652 7100
rect 2652 7044 2656 7100
rect 2592 7040 2656 7044
rect 7352 7100 7416 7104
rect 7352 7044 7356 7100
rect 7356 7044 7412 7100
rect 7412 7044 7416 7100
rect 7352 7040 7416 7044
rect 7432 7100 7496 7104
rect 7432 7044 7436 7100
rect 7436 7044 7492 7100
rect 7492 7044 7496 7100
rect 7432 7040 7496 7044
rect 7512 7100 7576 7104
rect 7512 7044 7516 7100
rect 7516 7044 7572 7100
rect 7572 7044 7576 7100
rect 7512 7040 7576 7044
rect 7592 7100 7656 7104
rect 7592 7044 7596 7100
rect 7596 7044 7652 7100
rect 7652 7044 7656 7100
rect 7592 7040 7656 7044
rect 6316 6836 6380 6900
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 8012 6556 8076 6560
rect 8012 6500 8016 6556
rect 8016 6500 8072 6556
rect 8072 6500 8076 6556
rect 8012 6496 8076 6500
rect 8092 6556 8156 6560
rect 8092 6500 8096 6556
rect 8096 6500 8152 6556
rect 8152 6500 8156 6556
rect 8092 6496 8156 6500
rect 8172 6556 8236 6560
rect 8172 6500 8176 6556
rect 8176 6500 8232 6556
rect 8232 6500 8236 6556
rect 8172 6496 8236 6500
rect 8252 6556 8316 6560
rect 8252 6500 8256 6556
rect 8256 6500 8312 6556
rect 8312 6500 8316 6556
rect 8252 6496 8316 6500
rect 2352 6012 2416 6016
rect 2352 5956 2356 6012
rect 2356 5956 2412 6012
rect 2412 5956 2416 6012
rect 2352 5952 2416 5956
rect 2432 6012 2496 6016
rect 2432 5956 2436 6012
rect 2436 5956 2492 6012
rect 2492 5956 2496 6012
rect 2432 5952 2496 5956
rect 2512 6012 2576 6016
rect 2512 5956 2516 6012
rect 2516 5956 2572 6012
rect 2572 5956 2576 6012
rect 2512 5952 2576 5956
rect 2592 6012 2656 6016
rect 2592 5956 2596 6012
rect 2596 5956 2652 6012
rect 2652 5956 2656 6012
rect 2592 5952 2656 5956
rect 7352 6012 7416 6016
rect 7352 5956 7356 6012
rect 7356 5956 7412 6012
rect 7412 5956 7416 6012
rect 7352 5952 7416 5956
rect 7432 6012 7496 6016
rect 7432 5956 7436 6012
rect 7436 5956 7492 6012
rect 7492 5956 7496 6012
rect 7432 5952 7496 5956
rect 7512 6012 7576 6016
rect 7512 5956 7516 6012
rect 7516 5956 7572 6012
rect 7572 5956 7576 6012
rect 7512 5952 7576 5956
rect 7592 6012 7656 6016
rect 7592 5956 7596 6012
rect 7596 5956 7652 6012
rect 7652 5956 7656 6012
rect 7592 5952 7656 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 8012 5468 8076 5472
rect 8012 5412 8016 5468
rect 8016 5412 8072 5468
rect 8072 5412 8076 5468
rect 8012 5408 8076 5412
rect 8092 5468 8156 5472
rect 8092 5412 8096 5468
rect 8096 5412 8152 5468
rect 8152 5412 8156 5468
rect 8092 5408 8156 5412
rect 8172 5468 8236 5472
rect 8172 5412 8176 5468
rect 8176 5412 8232 5468
rect 8232 5412 8236 5468
rect 8172 5408 8236 5412
rect 8252 5468 8316 5472
rect 8252 5412 8256 5468
rect 8256 5412 8312 5468
rect 8312 5412 8316 5468
rect 8252 5408 8316 5412
rect 2352 4924 2416 4928
rect 2352 4868 2356 4924
rect 2356 4868 2412 4924
rect 2412 4868 2416 4924
rect 2352 4864 2416 4868
rect 2432 4924 2496 4928
rect 2432 4868 2436 4924
rect 2436 4868 2492 4924
rect 2492 4868 2496 4924
rect 2432 4864 2496 4868
rect 2512 4924 2576 4928
rect 2512 4868 2516 4924
rect 2516 4868 2572 4924
rect 2572 4868 2576 4924
rect 2512 4864 2576 4868
rect 2592 4924 2656 4928
rect 2592 4868 2596 4924
rect 2596 4868 2652 4924
rect 2652 4868 2656 4924
rect 2592 4864 2656 4868
rect 7352 4924 7416 4928
rect 7352 4868 7356 4924
rect 7356 4868 7412 4924
rect 7412 4868 7416 4924
rect 7352 4864 7416 4868
rect 7432 4924 7496 4928
rect 7432 4868 7436 4924
rect 7436 4868 7492 4924
rect 7492 4868 7496 4924
rect 7432 4864 7496 4868
rect 7512 4924 7576 4928
rect 7512 4868 7516 4924
rect 7516 4868 7572 4924
rect 7572 4868 7576 4924
rect 7512 4864 7576 4868
rect 7592 4924 7656 4928
rect 7592 4868 7596 4924
rect 7596 4868 7652 4924
rect 7652 4868 7656 4924
rect 7592 4864 7656 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 8012 4380 8076 4384
rect 8012 4324 8016 4380
rect 8016 4324 8072 4380
rect 8072 4324 8076 4380
rect 8012 4320 8076 4324
rect 8092 4380 8156 4384
rect 8092 4324 8096 4380
rect 8096 4324 8152 4380
rect 8152 4324 8156 4380
rect 8092 4320 8156 4324
rect 8172 4380 8236 4384
rect 8172 4324 8176 4380
rect 8176 4324 8232 4380
rect 8232 4324 8236 4380
rect 8172 4320 8236 4324
rect 8252 4380 8316 4384
rect 8252 4324 8256 4380
rect 8256 4324 8312 4380
rect 8312 4324 8316 4380
rect 8252 4320 8316 4324
rect 2352 3836 2416 3840
rect 2352 3780 2356 3836
rect 2356 3780 2412 3836
rect 2412 3780 2416 3836
rect 2352 3776 2416 3780
rect 2432 3836 2496 3840
rect 2432 3780 2436 3836
rect 2436 3780 2492 3836
rect 2492 3780 2496 3836
rect 2432 3776 2496 3780
rect 2512 3836 2576 3840
rect 2512 3780 2516 3836
rect 2516 3780 2572 3836
rect 2572 3780 2576 3836
rect 2512 3776 2576 3780
rect 2592 3836 2656 3840
rect 2592 3780 2596 3836
rect 2596 3780 2652 3836
rect 2652 3780 2656 3836
rect 2592 3776 2656 3780
rect 7352 3836 7416 3840
rect 7352 3780 7356 3836
rect 7356 3780 7412 3836
rect 7412 3780 7416 3836
rect 7352 3776 7416 3780
rect 7432 3836 7496 3840
rect 7432 3780 7436 3836
rect 7436 3780 7492 3836
rect 7492 3780 7496 3836
rect 7432 3776 7496 3780
rect 7512 3836 7576 3840
rect 7512 3780 7516 3836
rect 7516 3780 7572 3836
rect 7572 3780 7576 3836
rect 7512 3776 7576 3780
rect 7592 3836 7656 3840
rect 7592 3780 7596 3836
rect 7596 3780 7652 3836
rect 7652 3780 7656 3836
rect 7592 3776 7656 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 8012 3292 8076 3296
rect 8012 3236 8016 3292
rect 8016 3236 8072 3292
rect 8072 3236 8076 3292
rect 8012 3232 8076 3236
rect 8092 3292 8156 3296
rect 8092 3236 8096 3292
rect 8096 3236 8152 3292
rect 8152 3236 8156 3292
rect 8092 3232 8156 3236
rect 8172 3292 8236 3296
rect 8172 3236 8176 3292
rect 8176 3236 8232 3292
rect 8232 3236 8236 3292
rect 8172 3232 8236 3236
rect 8252 3292 8316 3296
rect 8252 3236 8256 3292
rect 8256 3236 8312 3292
rect 8312 3236 8316 3292
rect 8252 3232 8316 3236
rect 2352 2748 2416 2752
rect 2352 2692 2356 2748
rect 2356 2692 2412 2748
rect 2412 2692 2416 2748
rect 2352 2688 2416 2692
rect 2432 2748 2496 2752
rect 2432 2692 2436 2748
rect 2436 2692 2492 2748
rect 2492 2692 2496 2748
rect 2432 2688 2496 2692
rect 2512 2748 2576 2752
rect 2512 2692 2516 2748
rect 2516 2692 2572 2748
rect 2572 2692 2576 2748
rect 2512 2688 2576 2692
rect 2592 2748 2656 2752
rect 2592 2692 2596 2748
rect 2596 2692 2652 2748
rect 2652 2692 2656 2748
rect 2592 2688 2656 2692
rect 7352 2748 7416 2752
rect 7352 2692 7356 2748
rect 7356 2692 7412 2748
rect 7412 2692 7416 2748
rect 7352 2688 7416 2692
rect 7432 2748 7496 2752
rect 7432 2692 7436 2748
rect 7436 2692 7492 2748
rect 7492 2692 7496 2748
rect 7432 2688 7496 2692
rect 7512 2748 7576 2752
rect 7512 2692 7516 2748
rect 7516 2692 7572 2748
rect 7572 2692 7576 2748
rect 7512 2688 7576 2692
rect 7592 2748 7656 2752
rect 7592 2692 7596 2748
rect 7596 2692 7652 2748
rect 7652 2692 7656 2748
rect 7592 2688 7656 2692
rect 6684 2680 6748 2684
rect 6684 2624 6698 2680
rect 6698 2624 6748 2680
rect 6684 2620 6748 2624
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 8012 2204 8076 2208
rect 8012 2148 8016 2204
rect 8016 2148 8072 2204
rect 8072 2148 8076 2204
rect 8012 2144 8076 2148
rect 8092 2204 8156 2208
rect 8092 2148 8096 2204
rect 8096 2148 8152 2204
rect 8152 2148 8156 2204
rect 8092 2144 8156 2148
rect 8172 2204 8236 2208
rect 8172 2148 8176 2204
rect 8176 2148 8232 2204
rect 8232 2148 8236 2204
rect 8172 2144 8236 2148
rect 8252 2204 8316 2208
rect 8252 2148 8256 2204
rect 8256 2148 8312 2204
rect 8312 2148 8316 2204
rect 8252 2144 8316 2148
<< metal4 >>
rect -1076 79930 -756 79972
rect -1076 79694 -1034 79930
rect -798 79694 -756 79930
rect -1076 74354 -756 79694
rect -1076 74118 -1034 74354
rect -798 74118 -756 74354
rect -1076 69354 -756 74118
rect -1076 69118 -1034 69354
rect -798 69118 -756 69354
rect -1076 64354 -756 69118
rect -1076 64118 -1034 64354
rect -798 64118 -756 64354
rect -1076 59354 -756 64118
rect -1076 59118 -1034 59354
rect -798 59118 -756 59354
rect -1076 54354 -756 59118
rect -1076 54118 -1034 54354
rect -798 54118 -756 54354
rect -1076 49354 -756 54118
rect -1076 49118 -1034 49354
rect -798 49118 -756 49354
rect -1076 44354 -756 49118
rect -1076 44118 -1034 44354
rect -798 44118 -756 44354
rect -1076 39354 -756 44118
rect -1076 39118 -1034 39354
rect -798 39118 -756 39354
rect -1076 34354 -756 39118
rect -1076 34118 -1034 34354
rect -798 34118 -756 34354
rect -1076 29354 -756 34118
rect -1076 29118 -1034 29354
rect -798 29118 -756 29354
rect -1076 24354 -756 29118
rect -1076 24118 -1034 24354
rect -798 24118 -756 24354
rect -1076 19354 -756 24118
rect -1076 19118 -1034 19354
rect -798 19118 -756 19354
rect -1076 14354 -756 19118
rect -1076 14118 -1034 14354
rect -798 14118 -756 14354
rect -1076 9354 -756 14118
rect -1076 9118 -1034 9354
rect -798 9118 -756 9354
rect -1076 4354 -756 9118
rect -1076 4118 -1034 4354
rect -798 4118 -756 4354
rect -1076 274 -756 4118
rect -416 79270 -96 79312
rect -416 79034 -374 79270
rect -138 79034 -96 79270
rect -416 73694 -96 79034
rect -416 73458 -374 73694
rect -138 73458 -96 73694
rect -416 68694 -96 73458
rect -416 68458 -374 68694
rect -138 68458 -96 68694
rect -416 63694 -96 68458
rect -416 63458 -374 63694
rect -138 63458 -96 63694
rect -416 58694 -96 63458
rect -416 58458 -374 58694
rect -138 58458 -96 58694
rect -416 53694 -96 58458
rect -416 53458 -374 53694
rect -138 53458 -96 53694
rect -416 48694 -96 53458
rect -416 48458 -374 48694
rect -138 48458 -96 48694
rect -416 43694 -96 48458
rect -416 43458 -374 43694
rect -138 43458 -96 43694
rect -416 38694 -96 43458
rect -416 38458 -374 38694
rect -138 38458 -96 38694
rect -416 33694 -96 38458
rect -416 33458 -374 33694
rect -138 33458 -96 33694
rect -416 28694 -96 33458
rect -416 28458 -374 28694
rect -138 28458 -96 28694
rect -416 23694 -96 28458
rect -416 23458 -374 23694
rect -138 23458 -96 23694
rect -416 18694 -96 23458
rect -416 18458 -374 18694
rect -138 18458 -96 18694
rect -416 13694 -96 18458
rect -416 13458 -374 13694
rect -138 13458 -96 13694
rect -416 8694 -96 13458
rect -416 8458 -374 8694
rect -138 8458 -96 8694
rect -416 3694 -96 8458
rect -416 3458 -374 3694
rect -138 3458 -96 3694
rect -416 934 -96 3458
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 2344 79270 2664 79972
rect 2344 79034 2386 79270
rect 2622 79034 2664 79270
rect 2344 77824 2664 79034
rect 2344 77760 2352 77824
rect 2416 77760 2432 77824
rect 2496 77760 2512 77824
rect 2576 77760 2592 77824
rect 2656 77760 2664 77824
rect 2344 76736 2664 77760
rect 2344 76672 2352 76736
rect 2416 76672 2432 76736
rect 2496 76672 2512 76736
rect 2576 76672 2592 76736
rect 2656 76672 2664 76736
rect 2344 75648 2664 76672
rect 2344 75584 2352 75648
rect 2416 75584 2432 75648
rect 2496 75584 2512 75648
rect 2576 75584 2592 75648
rect 2656 75584 2664 75648
rect 2344 74560 2664 75584
rect 2344 74496 2352 74560
rect 2416 74496 2432 74560
rect 2496 74496 2512 74560
rect 2576 74496 2592 74560
rect 2656 74496 2664 74560
rect 2344 73694 2664 74496
rect 2344 73472 2386 73694
rect 2622 73472 2664 73694
rect 2344 73408 2352 73472
rect 2416 73408 2432 73458
rect 2496 73408 2512 73458
rect 2576 73408 2592 73458
rect 2656 73408 2664 73472
rect 2344 72384 2664 73408
rect 2344 72320 2352 72384
rect 2416 72320 2432 72384
rect 2496 72320 2512 72384
rect 2576 72320 2592 72384
rect 2656 72320 2664 72384
rect 2344 71296 2664 72320
rect 2344 71232 2352 71296
rect 2416 71232 2432 71296
rect 2496 71232 2512 71296
rect 2576 71232 2592 71296
rect 2656 71232 2664 71296
rect 2344 70208 2664 71232
rect 2344 70144 2352 70208
rect 2416 70144 2432 70208
rect 2496 70144 2512 70208
rect 2576 70144 2592 70208
rect 2656 70144 2664 70208
rect 2344 69120 2664 70144
rect 2344 69056 2352 69120
rect 2416 69056 2432 69120
rect 2496 69056 2512 69120
rect 2576 69056 2592 69120
rect 2656 69056 2664 69120
rect 2344 68694 2664 69056
rect 2344 68458 2386 68694
rect 2622 68458 2664 68694
rect 2344 68032 2664 68458
rect 2344 67968 2352 68032
rect 2416 67968 2432 68032
rect 2496 67968 2512 68032
rect 2576 67968 2592 68032
rect 2656 67968 2664 68032
rect 2344 66944 2664 67968
rect 2344 66880 2352 66944
rect 2416 66880 2432 66944
rect 2496 66880 2512 66944
rect 2576 66880 2592 66944
rect 2656 66880 2664 66944
rect 2344 65856 2664 66880
rect 2344 65792 2352 65856
rect 2416 65792 2432 65856
rect 2496 65792 2512 65856
rect 2576 65792 2592 65856
rect 2656 65792 2664 65856
rect 2344 64768 2664 65792
rect 2344 64704 2352 64768
rect 2416 64704 2432 64768
rect 2496 64704 2512 64768
rect 2576 64704 2592 64768
rect 2656 64704 2664 64768
rect 2344 63694 2664 64704
rect 2344 63680 2386 63694
rect 2622 63680 2664 63694
rect 2344 63616 2352 63680
rect 2656 63616 2664 63680
rect 2344 63458 2386 63616
rect 2622 63458 2664 63616
rect 2344 62592 2664 63458
rect 2344 62528 2352 62592
rect 2416 62528 2432 62592
rect 2496 62528 2512 62592
rect 2576 62528 2592 62592
rect 2656 62528 2664 62592
rect 2344 61504 2664 62528
rect 2344 61440 2352 61504
rect 2416 61440 2432 61504
rect 2496 61440 2512 61504
rect 2576 61440 2592 61504
rect 2656 61440 2664 61504
rect 2344 60416 2664 61440
rect 2344 60352 2352 60416
rect 2416 60352 2432 60416
rect 2496 60352 2512 60416
rect 2576 60352 2592 60416
rect 2656 60352 2664 60416
rect 2344 59328 2664 60352
rect 2344 59264 2352 59328
rect 2416 59264 2432 59328
rect 2496 59264 2512 59328
rect 2576 59264 2592 59328
rect 2656 59264 2664 59328
rect 2344 58694 2664 59264
rect 2344 58458 2386 58694
rect 2622 58458 2664 58694
rect 2344 58240 2664 58458
rect 2344 58176 2352 58240
rect 2416 58176 2432 58240
rect 2496 58176 2512 58240
rect 2576 58176 2592 58240
rect 2656 58176 2664 58240
rect 2344 57152 2664 58176
rect 2344 57088 2352 57152
rect 2416 57088 2432 57152
rect 2496 57088 2512 57152
rect 2576 57088 2592 57152
rect 2656 57088 2664 57152
rect 2344 56064 2664 57088
rect 2344 56000 2352 56064
rect 2416 56000 2432 56064
rect 2496 56000 2512 56064
rect 2576 56000 2592 56064
rect 2656 56000 2664 56064
rect 2344 54976 2664 56000
rect 2344 54912 2352 54976
rect 2416 54912 2432 54976
rect 2496 54912 2512 54976
rect 2576 54912 2592 54976
rect 2656 54912 2664 54976
rect 2344 53888 2664 54912
rect 2344 53824 2352 53888
rect 2416 53824 2432 53888
rect 2496 53824 2512 53888
rect 2576 53824 2592 53888
rect 2656 53824 2664 53888
rect 2344 53694 2664 53824
rect 2344 53458 2386 53694
rect 2622 53458 2664 53694
rect 2344 52800 2664 53458
rect 2344 52736 2352 52800
rect 2416 52736 2432 52800
rect 2496 52736 2512 52800
rect 2576 52736 2592 52800
rect 2656 52736 2664 52800
rect 2344 51712 2664 52736
rect 2344 51648 2352 51712
rect 2416 51648 2432 51712
rect 2496 51648 2512 51712
rect 2576 51648 2592 51712
rect 2656 51648 2664 51712
rect 2344 50624 2664 51648
rect 2344 50560 2352 50624
rect 2416 50560 2432 50624
rect 2496 50560 2512 50624
rect 2576 50560 2592 50624
rect 2656 50560 2664 50624
rect 2344 49536 2664 50560
rect 2344 49472 2352 49536
rect 2416 49472 2432 49536
rect 2496 49472 2512 49536
rect 2576 49472 2592 49536
rect 2656 49472 2664 49536
rect 2344 48694 2664 49472
rect 2344 48458 2386 48694
rect 2622 48458 2664 48694
rect 2344 48448 2664 48458
rect 2344 48384 2352 48448
rect 2416 48384 2432 48448
rect 2496 48384 2512 48448
rect 2576 48384 2592 48448
rect 2656 48384 2664 48448
rect 2344 47360 2664 48384
rect 2344 47296 2352 47360
rect 2416 47296 2432 47360
rect 2496 47296 2512 47360
rect 2576 47296 2592 47360
rect 2656 47296 2664 47360
rect 2344 46272 2664 47296
rect 2344 46208 2352 46272
rect 2416 46208 2432 46272
rect 2496 46208 2512 46272
rect 2576 46208 2592 46272
rect 2656 46208 2664 46272
rect 2344 45184 2664 46208
rect 2344 45120 2352 45184
rect 2416 45120 2432 45184
rect 2496 45120 2512 45184
rect 2576 45120 2592 45184
rect 2656 45120 2664 45184
rect 2344 44096 2664 45120
rect 2344 44032 2352 44096
rect 2416 44032 2432 44096
rect 2496 44032 2512 44096
rect 2576 44032 2592 44096
rect 2656 44032 2664 44096
rect 2344 43694 2664 44032
rect 2344 43458 2386 43694
rect 2622 43458 2664 43694
rect 2344 43008 2664 43458
rect 2344 42944 2352 43008
rect 2416 42944 2432 43008
rect 2496 42944 2512 43008
rect 2576 42944 2592 43008
rect 2656 42944 2664 43008
rect 2344 41920 2664 42944
rect 2344 41856 2352 41920
rect 2416 41856 2432 41920
rect 2496 41856 2512 41920
rect 2576 41856 2592 41920
rect 2656 41856 2664 41920
rect 2344 40832 2664 41856
rect 2344 40768 2352 40832
rect 2416 40768 2432 40832
rect 2496 40768 2512 40832
rect 2576 40768 2592 40832
rect 2656 40768 2664 40832
rect 2344 39744 2664 40768
rect 2344 39680 2352 39744
rect 2416 39680 2432 39744
rect 2496 39680 2512 39744
rect 2576 39680 2592 39744
rect 2656 39680 2664 39744
rect 2344 38694 2664 39680
rect 2344 38656 2386 38694
rect 2622 38656 2664 38694
rect 2344 38592 2352 38656
rect 2656 38592 2664 38656
rect 2344 38458 2386 38592
rect 2622 38458 2664 38592
rect 2344 37568 2664 38458
rect 2344 37504 2352 37568
rect 2416 37504 2432 37568
rect 2496 37504 2512 37568
rect 2576 37504 2592 37568
rect 2656 37504 2664 37568
rect 2344 36480 2664 37504
rect 2344 36416 2352 36480
rect 2416 36416 2432 36480
rect 2496 36416 2512 36480
rect 2576 36416 2592 36480
rect 2656 36416 2664 36480
rect 2344 35392 2664 36416
rect 2344 35328 2352 35392
rect 2416 35328 2432 35392
rect 2496 35328 2512 35392
rect 2576 35328 2592 35392
rect 2656 35328 2664 35392
rect 2344 34304 2664 35328
rect 2344 34240 2352 34304
rect 2416 34240 2432 34304
rect 2496 34240 2512 34304
rect 2576 34240 2592 34304
rect 2656 34240 2664 34304
rect 2344 33694 2664 34240
rect 2344 33458 2386 33694
rect 2622 33458 2664 33694
rect 2344 33216 2664 33458
rect 2344 33152 2352 33216
rect 2416 33152 2432 33216
rect 2496 33152 2512 33216
rect 2576 33152 2592 33216
rect 2656 33152 2664 33216
rect 2344 32128 2664 33152
rect 2344 32064 2352 32128
rect 2416 32064 2432 32128
rect 2496 32064 2512 32128
rect 2576 32064 2592 32128
rect 2656 32064 2664 32128
rect 2344 31040 2664 32064
rect 2344 30976 2352 31040
rect 2416 30976 2432 31040
rect 2496 30976 2512 31040
rect 2576 30976 2592 31040
rect 2656 30976 2664 31040
rect 2344 29952 2664 30976
rect 2344 29888 2352 29952
rect 2416 29888 2432 29952
rect 2496 29888 2512 29952
rect 2576 29888 2592 29952
rect 2656 29888 2664 29952
rect 2344 28864 2664 29888
rect 2344 28800 2352 28864
rect 2416 28800 2432 28864
rect 2496 28800 2512 28864
rect 2576 28800 2592 28864
rect 2656 28800 2664 28864
rect 2344 28694 2664 28800
rect 2344 28458 2386 28694
rect 2622 28458 2664 28694
rect 2344 27776 2664 28458
rect 2344 27712 2352 27776
rect 2416 27712 2432 27776
rect 2496 27712 2512 27776
rect 2576 27712 2592 27776
rect 2656 27712 2664 27776
rect 2344 26688 2664 27712
rect 2344 26624 2352 26688
rect 2416 26624 2432 26688
rect 2496 26624 2512 26688
rect 2576 26624 2592 26688
rect 2656 26624 2664 26688
rect 2344 25600 2664 26624
rect 2344 25536 2352 25600
rect 2416 25536 2432 25600
rect 2496 25536 2512 25600
rect 2576 25536 2592 25600
rect 2656 25536 2664 25600
rect 2344 24512 2664 25536
rect 2344 24448 2352 24512
rect 2416 24448 2432 24512
rect 2496 24448 2512 24512
rect 2576 24448 2592 24512
rect 2656 24448 2664 24512
rect 2344 23694 2664 24448
rect 2344 23458 2386 23694
rect 2622 23458 2664 23694
rect 2344 23424 2664 23458
rect 2344 23360 2352 23424
rect 2416 23360 2432 23424
rect 2496 23360 2512 23424
rect 2576 23360 2592 23424
rect 2656 23360 2664 23424
rect 2344 22336 2664 23360
rect 2344 22272 2352 22336
rect 2416 22272 2432 22336
rect 2496 22272 2512 22336
rect 2576 22272 2592 22336
rect 2656 22272 2664 22336
rect 2344 21248 2664 22272
rect 2344 21184 2352 21248
rect 2416 21184 2432 21248
rect 2496 21184 2512 21248
rect 2576 21184 2592 21248
rect 2656 21184 2664 21248
rect 2344 20160 2664 21184
rect 2344 20096 2352 20160
rect 2416 20096 2432 20160
rect 2496 20096 2512 20160
rect 2576 20096 2592 20160
rect 2656 20096 2664 20160
rect 2344 19072 2664 20096
rect 2344 19008 2352 19072
rect 2416 19008 2432 19072
rect 2496 19008 2512 19072
rect 2576 19008 2592 19072
rect 2656 19008 2664 19072
rect 2344 18694 2664 19008
rect 2344 18458 2386 18694
rect 2622 18458 2664 18694
rect 2344 17984 2664 18458
rect 2344 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2664 17984
rect 2344 16896 2664 17920
rect 2344 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2664 16896
rect 2344 15808 2664 16832
rect 2344 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2664 15808
rect 2344 14720 2664 15744
rect 2344 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2664 14720
rect 2344 13694 2664 14656
rect 2344 13632 2386 13694
rect 2622 13632 2664 13694
rect 2344 13568 2352 13632
rect 2656 13568 2664 13632
rect 2344 13458 2386 13568
rect 2622 13458 2664 13568
rect 2344 12544 2664 13458
rect 2344 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2664 12544
rect 2344 11456 2664 12480
rect 2344 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2664 11456
rect 2344 10368 2664 11392
rect 2344 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2664 10368
rect 2344 9280 2664 10304
rect 2344 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2664 9280
rect 2344 8694 2664 9216
rect 2344 8458 2386 8694
rect 2622 8458 2664 8694
rect 2344 8192 2664 8458
rect 2344 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2664 8192
rect 2344 7104 2664 8128
rect 2344 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2664 7104
rect 2344 6016 2664 7040
rect 2344 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2664 6016
rect 2344 4928 2664 5952
rect 2344 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2664 4928
rect 2344 3840 2664 4864
rect 2344 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2664 3840
rect 2344 3694 2664 3776
rect 2344 3458 2386 3694
rect 2622 3458 2664 3694
rect 2344 2752 2664 3458
rect 2344 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2664 2752
rect 2344 934 2664 2688
rect 2344 698 2386 934
rect 2622 698 2664 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 2344 -4 2664 698
rect 3004 79930 3324 79972
rect 3004 79694 3046 79930
rect 3282 79694 3324 79930
rect 3004 77280 3324 79694
rect 3004 77216 3012 77280
rect 3076 77216 3092 77280
rect 3156 77216 3172 77280
rect 3236 77216 3252 77280
rect 3316 77216 3324 77280
rect 3004 76192 3324 77216
rect 3004 76128 3012 76192
rect 3076 76128 3092 76192
rect 3156 76128 3172 76192
rect 3236 76128 3252 76192
rect 3316 76128 3324 76192
rect 3004 75104 3324 76128
rect 3004 75040 3012 75104
rect 3076 75040 3092 75104
rect 3156 75040 3172 75104
rect 3236 75040 3252 75104
rect 3316 75040 3324 75104
rect 3004 74354 3324 75040
rect 3004 74118 3046 74354
rect 3282 74118 3324 74354
rect 3004 74016 3324 74118
rect 3004 73952 3012 74016
rect 3076 73952 3092 74016
rect 3156 73952 3172 74016
rect 3236 73952 3252 74016
rect 3316 73952 3324 74016
rect 3004 72928 3324 73952
rect 3004 72864 3012 72928
rect 3076 72864 3092 72928
rect 3156 72864 3172 72928
rect 3236 72864 3252 72928
rect 3316 72864 3324 72928
rect 3004 71840 3324 72864
rect 3004 71776 3012 71840
rect 3076 71776 3092 71840
rect 3156 71776 3172 71840
rect 3236 71776 3252 71840
rect 3316 71776 3324 71840
rect 3004 70752 3324 71776
rect 3004 70688 3012 70752
rect 3076 70688 3092 70752
rect 3156 70688 3172 70752
rect 3236 70688 3252 70752
rect 3316 70688 3324 70752
rect 3004 69664 3324 70688
rect 3004 69600 3012 69664
rect 3076 69600 3092 69664
rect 3156 69600 3172 69664
rect 3236 69600 3252 69664
rect 3316 69600 3324 69664
rect 3004 69354 3324 69600
rect 3004 69118 3046 69354
rect 3282 69118 3324 69354
rect 3004 68576 3324 69118
rect 3004 68512 3012 68576
rect 3076 68512 3092 68576
rect 3156 68512 3172 68576
rect 3236 68512 3252 68576
rect 3316 68512 3324 68576
rect 3004 67488 3324 68512
rect 3004 67424 3012 67488
rect 3076 67424 3092 67488
rect 3156 67424 3172 67488
rect 3236 67424 3252 67488
rect 3316 67424 3324 67488
rect 3004 66400 3324 67424
rect 3004 66336 3012 66400
rect 3076 66336 3092 66400
rect 3156 66336 3172 66400
rect 3236 66336 3252 66400
rect 3316 66336 3324 66400
rect 3004 65312 3324 66336
rect 3004 65248 3012 65312
rect 3076 65248 3092 65312
rect 3156 65248 3172 65312
rect 3236 65248 3252 65312
rect 3316 65248 3324 65312
rect 3004 64354 3324 65248
rect 3004 64224 3046 64354
rect 3282 64224 3324 64354
rect 3004 64160 3012 64224
rect 3316 64160 3324 64224
rect 3004 64118 3046 64160
rect 3282 64118 3324 64160
rect 3004 63136 3324 64118
rect 3004 63072 3012 63136
rect 3076 63072 3092 63136
rect 3156 63072 3172 63136
rect 3236 63072 3252 63136
rect 3316 63072 3324 63136
rect 3004 62048 3324 63072
rect 3004 61984 3012 62048
rect 3076 61984 3092 62048
rect 3156 61984 3172 62048
rect 3236 61984 3252 62048
rect 3316 61984 3324 62048
rect 3004 60960 3324 61984
rect 3004 60896 3012 60960
rect 3076 60896 3092 60960
rect 3156 60896 3172 60960
rect 3236 60896 3252 60960
rect 3316 60896 3324 60960
rect 3004 59872 3324 60896
rect 3004 59808 3012 59872
rect 3076 59808 3092 59872
rect 3156 59808 3172 59872
rect 3236 59808 3252 59872
rect 3316 59808 3324 59872
rect 3004 59354 3324 59808
rect 3004 59118 3046 59354
rect 3282 59118 3324 59354
rect 3004 58784 3324 59118
rect 3004 58720 3012 58784
rect 3076 58720 3092 58784
rect 3156 58720 3172 58784
rect 3236 58720 3252 58784
rect 3316 58720 3324 58784
rect 3004 57696 3324 58720
rect 3004 57632 3012 57696
rect 3076 57632 3092 57696
rect 3156 57632 3172 57696
rect 3236 57632 3252 57696
rect 3316 57632 3324 57696
rect 3004 56608 3324 57632
rect 3004 56544 3012 56608
rect 3076 56544 3092 56608
rect 3156 56544 3172 56608
rect 3236 56544 3252 56608
rect 3316 56544 3324 56608
rect 3004 55520 3324 56544
rect 3004 55456 3012 55520
rect 3076 55456 3092 55520
rect 3156 55456 3172 55520
rect 3236 55456 3252 55520
rect 3316 55456 3324 55520
rect 3004 54432 3324 55456
rect 3004 54368 3012 54432
rect 3076 54368 3092 54432
rect 3156 54368 3172 54432
rect 3236 54368 3252 54432
rect 3316 54368 3324 54432
rect 3004 54354 3324 54368
rect 3004 54118 3046 54354
rect 3282 54118 3324 54354
rect 3004 53344 3324 54118
rect 3004 53280 3012 53344
rect 3076 53280 3092 53344
rect 3156 53280 3172 53344
rect 3236 53280 3252 53344
rect 3316 53280 3324 53344
rect 3004 52256 3324 53280
rect 3004 52192 3012 52256
rect 3076 52192 3092 52256
rect 3156 52192 3172 52256
rect 3236 52192 3252 52256
rect 3316 52192 3324 52256
rect 3004 51168 3324 52192
rect 3004 51104 3012 51168
rect 3076 51104 3092 51168
rect 3156 51104 3172 51168
rect 3236 51104 3252 51168
rect 3316 51104 3324 51168
rect 3004 50080 3324 51104
rect 3004 50016 3012 50080
rect 3076 50016 3092 50080
rect 3156 50016 3172 50080
rect 3236 50016 3252 50080
rect 3316 50016 3324 50080
rect 3004 49354 3324 50016
rect 3004 49118 3046 49354
rect 3282 49118 3324 49354
rect 3004 48992 3324 49118
rect 3004 48928 3012 48992
rect 3076 48928 3092 48992
rect 3156 48928 3172 48992
rect 3236 48928 3252 48992
rect 3316 48928 3324 48992
rect 3004 47904 3324 48928
rect 3004 47840 3012 47904
rect 3076 47840 3092 47904
rect 3156 47840 3172 47904
rect 3236 47840 3252 47904
rect 3316 47840 3324 47904
rect 3004 46816 3324 47840
rect 3004 46752 3012 46816
rect 3076 46752 3092 46816
rect 3156 46752 3172 46816
rect 3236 46752 3252 46816
rect 3316 46752 3324 46816
rect 3004 45728 3324 46752
rect 3004 45664 3012 45728
rect 3076 45664 3092 45728
rect 3156 45664 3172 45728
rect 3236 45664 3252 45728
rect 3316 45664 3324 45728
rect 3004 44640 3324 45664
rect 3004 44576 3012 44640
rect 3076 44576 3092 44640
rect 3156 44576 3172 44640
rect 3236 44576 3252 44640
rect 3316 44576 3324 44640
rect 3004 44354 3324 44576
rect 3004 44118 3046 44354
rect 3282 44118 3324 44354
rect 3004 43552 3324 44118
rect 3004 43488 3012 43552
rect 3076 43488 3092 43552
rect 3156 43488 3172 43552
rect 3236 43488 3252 43552
rect 3316 43488 3324 43552
rect 3004 42464 3324 43488
rect 3004 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3324 42464
rect 3004 41376 3324 42400
rect 7344 79270 7664 79972
rect 7344 79034 7386 79270
rect 7622 79034 7664 79270
rect 7344 77824 7664 79034
rect 7344 77760 7352 77824
rect 7416 77760 7432 77824
rect 7496 77760 7512 77824
rect 7576 77760 7592 77824
rect 7656 77760 7664 77824
rect 7344 76736 7664 77760
rect 7344 76672 7352 76736
rect 7416 76672 7432 76736
rect 7496 76672 7512 76736
rect 7576 76672 7592 76736
rect 7656 76672 7664 76736
rect 7344 75648 7664 76672
rect 7344 75584 7352 75648
rect 7416 75584 7432 75648
rect 7496 75584 7512 75648
rect 7576 75584 7592 75648
rect 7656 75584 7664 75648
rect 7344 74560 7664 75584
rect 7344 74496 7352 74560
rect 7416 74496 7432 74560
rect 7496 74496 7512 74560
rect 7576 74496 7592 74560
rect 7656 74496 7664 74560
rect 7344 73694 7664 74496
rect 7344 73472 7386 73694
rect 7622 73472 7664 73694
rect 7344 73408 7352 73472
rect 7416 73408 7432 73458
rect 7496 73408 7512 73458
rect 7576 73408 7592 73458
rect 7656 73408 7664 73472
rect 7344 72384 7664 73408
rect 7344 72320 7352 72384
rect 7416 72320 7432 72384
rect 7496 72320 7512 72384
rect 7576 72320 7592 72384
rect 7656 72320 7664 72384
rect 7344 71296 7664 72320
rect 7344 71232 7352 71296
rect 7416 71232 7432 71296
rect 7496 71232 7512 71296
rect 7576 71232 7592 71296
rect 7656 71232 7664 71296
rect 7344 70208 7664 71232
rect 7344 70144 7352 70208
rect 7416 70144 7432 70208
rect 7496 70144 7512 70208
rect 7576 70144 7592 70208
rect 7656 70144 7664 70208
rect 7344 69120 7664 70144
rect 7344 69056 7352 69120
rect 7416 69056 7432 69120
rect 7496 69056 7512 69120
rect 7576 69056 7592 69120
rect 7656 69056 7664 69120
rect 7344 68694 7664 69056
rect 7344 68458 7386 68694
rect 7622 68458 7664 68694
rect 7344 68032 7664 68458
rect 7344 67968 7352 68032
rect 7416 67968 7432 68032
rect 7496 67968 7512 68032
rect 7576 67968 7592 68032
rect 7656 67968 7664 68032
rect 7344 66944 7664 67968
rect 7344 66880 7352 66944
rect 7416 66880 7432 66944
rect 7496 66880 7512 66944
rect 7576 66880 7592 66944
rect 7656 66880 7664 66944
rect 7344 65856 7664 66880
rect 7344 65792 7352 65856
rect 7416 65792 7432 65856
rect 7496 65792 7512 65856
rect 7576 65792 7592 65856
rect 7656 65792 7664 65856
rect 7344 64768 7664 65792
rect 7344 64704 7352 64768
rect 7416 64704 7432 64768
rect 7496 64704 7512 64768
rect 7576 64704 7592 64768
rect 7656 64704 7664 64768
rect 7344 63694 7664 64704
rect 7344 63680 7386 63694
rect 7622 63680 7664 63694
rect 7344 63616 7352 63680
rect 7656 63616 7664 63680
rect 7344 63458 7386 63616
rect 7622 63458 7664 63616
rect 7344 62592 7664 63458
rect 7344 62528 7352 62592
rect 7416 62528 7432 62592
rect 7496 62528 7512 62592
rect 7576 62528 7592 62592
rect 7656 62528 7664 62592
rect 7344 61504 7664 62528
rect 7344 61440 7352 61504
rect 7416 61440 7432 61504
rect 7496 61440 7512 61504
rect 7576 61440 7592 61504
rect 7656 61440 7664 61504
rect 7344 60416 7664 61440
rect 7344 60352 7352 60416
rect 7416 60352 7432 60416
rect 7496 60352 7512 60416
rect 7576 60352 7592 60416
rect 7656 60352 7664 60416
rect 7344 59328 7664 60352
rect 7344 59264 7352 59328
rect 7416 59264 7432 59328
rect 7496 59264 7512 59328
rect 7576 59264 7592 59328
rect 7656 59264 7664 59328
rect 7344 58694 7664 59264
rect 7344 58458 7386 58694
rect 7622 58458 7664 58694
rect 7344 58240 7664 58458
rect 7344 58176 7352 58240
rect 7416 58176 7432 58240
rect 7496 58176 7512 58240
rect 7576 58176 7592 58240
rect 7656 58176 7664 58240
rect 7344 57152 7664 58176
rect 7344 57088 7352 57152
rect 7416 57088 7432 57152
rect 7496 57088 7512 57152
rect 7576 57088 7592 57152
rect 7656 57088 7664 57152
rect 7344 56064 7664 57088
rect 7344 56000 7352 56064
rect 7416 56000 7432 56064
rect 7496 56000 7512 56064
rect 7576 56000 7592 56064
rect 7656 56000 7664 56064
rect 7344 54976 7664 56000
rect 7344 54912 7352 54976
rect 7416 54912 7432 54976
rect 7496 54912 7512 54976
rect 7576 54912 7592 54976
rect 7656 54912 7664 54976
rect 7344 53888 7664 54912
rect 7344 53824 7352 53888
rect 7416 53824 7432 53888
rect 7496 53824 7512 53888
rect 7576 53824 7592 53888
rect 7656 53824 7664 53888
rect 7344 53694 7664 53824
rect 7344 53458 7386 53694
rect 7622 53458 7664 53694
rect 7344 52800 7664 53458
rect 7344 52736 7352 52800
rect 7416 52736 7432 52800
rect 7496 52736 7512 52800
rect 7576 52736 7592 52800
rect 7656 52736 7664 52800
rect 7344 51712 7664 52736
rect 7344 51648 7352 51712
rect 7416 51648 7432 51712
rect 7496 51648 7512 51712
rect 7576 51648 7592 51712
rect 7656 51648 7664 51712
rect 7344 50624 7664 51648
rect 7344 50560 7352 50624
rect 7416 50560 7432 50624
rect 7496 50560 7512 50624
rect 7576 50560 7592 50624
rect 7656 50560 7664 50624
rect 7344 49536 7664 50560
rect 7344 49472 7352 49536
rect 7416 49472 7432 49536
rect 7496 49472 7512 49536
rect 7576 49472 7592 49536
rect 7656 49472 7664 49536
rect 7344 48694 7664 49472
rect 7344 48458 7386 48694
rect 7622 48458 7664 48694
rect 7344 48448 7664 48458
rect 7344 48384 7352 48448
rect 7416 48384 7432 48448
rect 7496 48384 7512 48448
rect 7576 48384 7592 48448
rect 7656 48384 7664 48448
rect 7344 47360 7664 48384
rect 7344 47296 7352 47360
rect 7416 47296 7432 47360
rect 7496 47296 7512 47360
rect 7576 47296 7592 47360
rect 7656 47296 7664 47360
rect 7344 46272 7664 47296
rect 7344 46208 7352 46272
rect 7416 46208 7432 46272
rect 7496 46208 7512 46272
rect 7576 46208 7592 46272
rect 7656 46208 7664 46272
rect 7344 45184 7664 46208
rect 7344 45120 7352 45184
rect 7416 45120 7432 45184
rect 7496 45120 7512 45184
rect 7576 45120 7592 45184
rect 7656 45120 7664 45184
rect 7344 44096 7664 45120
rect 7344 44032 7352 44096
rect 7416 44032 7432 44096
rect 7496 44032 7512 44096
rect 7576 44032 7592 44096
rect 7656 44032 7664 44096
rect 7344 43694 7664 44032
rect 7344 43458 7386 43694
rect 7622 43458 7664 43694
rect 7344 43008 7664 43458
rect 7344 42944 7352 43008
rect 7416 42944 7432 43008
rect 7496 42944 7512 43008
rect 7576 42944 7592 43008
rect 7656 42944 7664 43008
rect 7344 41920 7664 42944
rect 7344 41856 7352 41920
rect 7416 41856 7432 41920
rect 7496 41856 7512 41920
rect 7576 41856 7592 41920
rect 7656 41856 7664 41920
rect 6315 41444 6381 41445
rect 6315 41380 6316 41444
rect 6380 41380 6381 41444
rect 6315 41379 6381 41380
rect 3004 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3324 41376
rect 3004 40288 3324 41312
rect 3004 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3324 40288
rect 3004 39354 3324 40224
rect 3004 39200 3046 39354
rect 3282 39200 3324 39354
rect 3004 39136 3012 39200
rect 3316 39136 3324 39200
rect 3004 39118 3046 39136
rect 3282 39118 3324 39136
rect 3004 38112 3324 39118
rect 3004 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3324 38112
rect 3004 37024 3324 38048
rect 3004 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3324 37024
rect 3004 35936 3324 36960
rect 3004 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3324 35936
rect 3004 34848 3324 35872
rect 3004 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3324 34848
rect 3004 34354 3324 34784
rect 3004 34118 3046 34354
rect 3282 34118 3324 34354
rect 3004 33760 3324 34118
rect 3004 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3324 33760
rect 3004 32672 3324 33696
rect 3004 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3324 32672
rect 3004 31584 3324 32608
rect 3004 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3324 31584
rect 3004 30496 3324 31520
rect 3004 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3324 30496
rect 3004 29408 3324 30432
rect 3004 29344 3012 29408
rect 3076 29354 3092 29408
rect 3156 29354 3172 29408
rect 3236 29354 3252 29408
rect 3316 29344 3324 29408
rect 3004 29118 3046 29344
rect 3282 29118 3324 29344
rect 3004 28320 3324 29118
rect 3004 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3324 28320
rect 3004 27232 3324 28256
rect 3004 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3324 27232
rect 3004 26144 3324 27168
rect 3004 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3324 26144
rect 3004 25056 3324 26080
rect 3004 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3324 25056
rect 3004 24354 3324 24992
rect 3004 24118 3046 24354
rect 3282 24118 3324 24354
rect 3004 23968 3324 24118
rect 3004 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3324 23968
rect 3004 22880 3324 23904
rect 3004 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3324 22880
rect 3004 21792 3324 22816
rect 3004 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3324 21792
rect 3004 20704 3324 21728
rect 3004 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3324 20704
rect 3004 19616 3324 20640
rect 3004 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3324 19616
rect 3004 19354 3324 19552
rect 3004 19118 3046 19354
rect 3282 19118 3324 19354
rect 3004 18528 3324 19118
rect 3004 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3324 18528
rect 3004 17440 3324 18464
rect 3004 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3324 17440
rect 3004 16352 3324 17376
rect 3004 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3324 16352
rect 3004 15264 3324 16288
rect 3004 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3324 15264
rect 3004 14354 3324 15200
rect 3004 14176 3046 14354
rect 3282 14176 3324 14354
rect 3004 14112 3012 14176
rect 3076 14112 3092 14118
rect 3156 14112 3172 14118
rect 3236 14112 3252 14118
rect 3316 14112 3324 14176
rect 3004 13088 3324 14112
rect 3004 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3324 13088
rect 3004 12000 3324 13024
rect 3004 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3324 12000
rect 3004 10912 3324 11936
rect 3004 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3324 10912
rect 3004 9824 3324 10848
rect 3004 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3324 9824
rect 3004 9354 3324 9760
rect 3004 9118 3046 9354
rect 3282 9118 3324 9354
rect 3004 8736 3324 9118
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 6318 6901 6378 41379
rect 7344 40832 7664 41856
rect 7344 40768 7352 40832
rect 7416 40768 7432 40832
rect 7496 40768 7512 40832
rect 7576 40768 7592 40832
rect 7656 40768 7664 40832
rect 6683 40084 6749 40085
rect 6683 40020 6684 40084
rect 6748 40020 6749 40084
rect 6683 40019 6749 40020
rect 6315 6900 6381 6901
rect 6315 6836 6316 6900
rect 6380 6836 6381 6900
rect 6315 6835 6381 6836
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4354 3092 4384
rect 3156 4354 3172 4384
rect 3236 4354 3252 4384
rect 3316 4320 3324 4384
rect 3004 4118 3046 4320
rect 3282 4118 3324 4320
rect 3004 3296 3324 4118
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 6686 2685 6746 40019
rect 7344 39744 7664 40768
rect 7344 39680 7352 39744
rect 7416 39680 7432 39744
rect 7496 39680 7512 39744
rect 7576 39680 7592 39744
rect 7656 39680 7664 39744
rect 7344 38694 7664 39680
rect 7344 38656 7386 38694
rect 7622 38656 7664 38694
rect 7344 38592 7352 38656
rect 7656 38592 7664 38656
rect 7344 38458 7386 38592
rect 7622 38458 7664 38592
rect 7344 37568 7664 38458
rect 7344 37504 7352 37568
rect 7416 37504 7432 37568
rect 7496 37504 7512 37568
rect 7576 37504 7592 37568
rect 7656 37504 7664 37568
rect 7344 36480 7664 37504
rect 7344 36416 7352 36480
rect 7416 36416 7432 36480
rect 7496 36416 7512 36480
rect 7576 36416 7592 36480
rect 7656 36416 7664 36480
rect 7344 35392 7664 36416
rect 7344 35328 7352 35392
rect 7416 35328 7432 35392
rect 7496 35328 7512 35392
rect 7576 35328 7592 35392
rect 7656 35328 7664 35392
rect 7344 34304 7664 35328
rect 7344 34240 7352 34304
rect 7416 34240 7432 34304
rect 7496 34240 7512 34304
rect 7576 34240 7592 34304
rect 7656 34240 7664 34304
rect 7344 33694 7664 34240
rect 7344 33458 7386 33694
rect 7622 33458 7664 33694
rect 7344 33216 7664 33458
rect 7344 33152 7352 33216
rect 7416 33152 7432 33216
rect 7496 33152 7512 33216
rect 7576 33152 7592 33216
rect 7656 33152 7664 33216
rect 7344 32128 7664 33152
rect 7344 32064 7352 32128
rect 7416 32064 7432 32128
rect 7496 32064 7512 32128
rect 7576 32064 7592 32128
rect 7656 32064 7664 32128
rect 7344 31040 7664 32064
rect 7344 30976 7352 31040
rect 7416 30976 7432 31040
rect 7496 30976 7512 31040
rect 7576 30976 7592 31040
rect 7656 30976 7664 31040
rect 7344 29952 7664 30976
rect 7344 29888 7352 29952
rect 7416 29888 7432 29952
rect 7496 29888 7512 29952
rect 7576 29888 7592 29952
rect 7656 29888 7664 29952
rect 7344 28864 7664 29888
rect 7344 28800 7352 28864
rect 7416 28800 7432 28864
rect 7496 28800 7512 28864
rect 7576 28800 7592 28864
rect 7656 28800 7664 28864
rect 7344 28694 7664 28800
rect 7344 28458 7386 28694
rect 7622 28458 7664 28694
rect 7344 27776 7664 28458
rect 7344 27712 7352 27776
rect 7416 27712 7432 27776
rect 7496 27712 7512 27776
rect 7576 27712 7592 27776
rect 7656 27712 7664 27776
rect 7344 26688 7664 27712
rect 7344 26624 7352 26688
rect 7416 26624 7432 26688
rect 7496 26624 7512 26688
rect 7576 26624 7592 26688
rect 7656 26624 7664 26688
rect 7344 25600 7664 26624
rect 7344 25536 7352 25600
rect 7416 25536 7432 25600
rect 7496 25536 7512 25600
rect 7576 25536 7592 25600
rect 7656 25536 7664 25600
rect 7344 24512 7664 25536
rect 7344 24448 7352 24512
rect 7416 24448 7432 24512
rect 7496 24448 7512 24512
rect 7576 24448 7592 24512
rect 7656 24448 7664 24512
rect 7344 23694 7664 24448
rect 7344 23458 7386 23694
rect 7622 23458 7664 23694
rect 7344 23424 7664 23458
rect 7344 23360 7352 23424
rect 7416 23360 7432 23424
rect 7496 23360 7512 23424
rect 7576 23360 7592 23424
rect 7656 23360 7664 23424
rect 7344 22336 7664 23360
rect 7344 22272 7352 22336
rect 7416 22272 7432 22336
rect 7496 22272 7512 22336
rect 7576 22272 7592 22336
rect 7656 22272 7664 22336
rect 7344 21248 7664 22272
rect 7344 21184 7352 21248
rect 7416 21184 7432 21248
rect 7496 21184 7512 21248
rect 7576 21184 7592 21248
rect 7656 21184 7664 21248
rect 7344 20160 7664 21184
rect 7344 20096 7352 20160
rect 7416 20096 7432 20160
rect 7496 20096 7512 20160
rect 7576 20096 7592 20160
rect 7656 20096 7664 20160
rect 7344 19072 7664 20096
rect 7344 19008 7352 19072
rect 7416 19008 7432 19072
rect 7496 19008 7512 19072
rect 7576 19008 7592 19072
rect 7656 19008 7664 19072
rect 7344 18694 7664 19008
rect 7344 18458 7386 18694
rect 7622 18458 7664 18694
rect 7344 17984 7664 18458
rect 7344 17920 7352 17984
rect 7416 17920 7432 17984
rect 7496 17920 7512 17984
rect 7576 17920 7592 17984
rect 7656 17920 7664 17984
rect 7344 16896 7664 17920
rect 7344 16832 7352 16896
rect 7416 16832 7432 16896
rect 7496 16832 7512 16896
rect 7576 16832 7592 16896
rect 7656 16832 7664 16896
rect 7344 15808 7664 16832
rect 7344 15744 7352 15808
rect 7416 15744 7432 15808
rect 7496 15744 7512 15808
rect 7576 15744 7592 15808
rect 7656 15744 7664 15808
rect 7344 14720 7664 15744
rect 7344 14656 7352 14720
rect 7416 14656 7432 14720
rect 7496 14656 7512 14720
rect 7576 14656 7592 14720
rect 7656 14656 7664 14720
rect 7344 13694 7664 14656
rect 7344 13632 7386 13694
rect 7622 13632 7664 13694
rect 7344 13568 7352 13632
rect 7656 13568 7664 13632
rect 7344 13458 7386 13568
rect 7622 13458 7664 13568
rect 7344 12544 7664 13458
rect 7344 12480 7352 12544
rect 7416 12480 7432 12544
rect 7496 12480 7512 12544
rect 7576 12480 7592 12544
rect 7656 12480 7664 12544
rect 7344 11456 7664 12480
rect 7344 11392 7352 11456
rect 7416 11392 7432 11456
rect 7496 11392 7512 11456
rect 7576 11392 7592 11456
rect 7656 11392 7664 11456
rect 7344 10368 7664 11392
rect 7344 10304 7352 10368
rect 7416 10304 7432 10368
rect 7496 10304 7512 10368
rect 7576 10304 7592 10368
rect 7656 10304 7664 10368
rect 7344 9280 7664 10304
rect 7344 9216 7352 9280
rect 7416 9216 7432 9280
rect 7496 9216 7512 9280
rect 7576 9216 7592 9280
rect 7656 9216 7664 9280
rect 7344 8694 7664 9216
rect 7344 8458 7386 8694
rect 7622 8458 7664 8694
rect 7344 8192 7664 8458
rect 7344 8128 7352 8192
rect 7416 8128 7432 8192
rect 7496 8128 7512 8192
rect 7576 8128 7592 8192
rect 7656 8128 7664 8192
rect 7344 7104 7664 8128
rect 7344 7040 7352 7104
rect 7416 7040 7432 7104
rect 7496 7040 7512 7104
rect 7576 7040 7592 7104
rect 7656 7040 7664 7104
rect 7344 6016 7664 7040
rect 7344 5952 7352 6016
rect 7416 5952 7432 6016
rect 7496 5952 7512 6016
rect 7576 5952 7592 6016
rect 7656 5952 7664 6016
rect 7344 4928 7664 5952
rect 7344 4864 7352 4928
rect 7416 4864 7432 4928
rect 7496 4864 7512 4928
rect 7576 4864 7592 4928
rect 7656 4864 7664 4928
rect 7344 3840 7664 4864
rect 7344 3776 7352 3840
rect 7416 3776 7432 3840
rect 7496 3776 7512 3840
rect 7576 3776 7592 3840
rect 7656 3776 7664 3840
rect 7344 3694 7664 3776
rect 7344 3458 7386 3694
rect 7622 3458 7664 3694
rect 7344 2752 7664 3458
rect 7344 2688 7352 2752
rect 7416 2688 7432 2752
rect 7496 2688 7512 2752
rect 7576 2688 7592 2752
rect 7656 2688 7664 2752
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 274 3324 2144
rect 3004 38 3046 274
rect 3282 38 3324 274
rect 3004 -4 3324 38
rect 7344 934 7664 2688
rect 7344 698 7386 934
rect 7622 698 7664 934
rect 7344 -4 7664 698
rect 8004 79930 8324 79972
rect 8004 79694 8046 79930
rect 8282 79694 8324 79930
rect 8004 77280 8324 79694
rect 10692 79930 11012 79972
rect 10692 79694 10734 79930
rect 10970 79694 11012 79930
rect 8004 77216 8012 77280
rect 8076 77216 8092 77280
rect 8156 77216 8172 77280
rect 8236 77216 8252 77280
rect 8316 77216 8324 77280
rect 8004 76192 8324 77216
rect 8004 76128 8012 76192
rect 8076 76128 8092 76192
rect 8156 76128 8172 76192
rect 8236 76128 8252 76192
rect 8316 76128 8324 76192
rect 8004 75104 8324 76128
rect 8004 75040 8012 75104
rect 8076 75040 8092 75104
rect 8156 75040 8172 75104
rect 8236 75040 8252 75104
rect 8316 75040 8324 75104
rect 8004 74354 8324 75040
rect 8004 74118 8046 74354
rect 8282 74118 8324 74354
rect 8004 74016 8324 74118
rect 8004 73952 8012 74016
rect 8076 73952 8092 74016
rect 8156 73952 8172 74016
rect 8236 73952 8252 74016
rect 8316 73952 8324 74016
rect 8004 72928 8324 73952
rect 8004 72864 8012 72928
rect 8076 72864 8092 72928
rect 8156 72864 8172 72928
rect 8236 72864 8252 72928
rect 8316 72864 8324 72928
rect 8004 71840 8324 72864
rect 8004 71776 8012 71840
rect 8076 71776 8092 71840
rect 8156 71776 8172 71840
rect 8236 71776 8252 71840
rect 8316 71776 8324 71840
rect 8004 70752 8324 71776
rect 8004 70688 8012 70752
rect 8076 70688 8092 70752
rect 8156 70688 8172 70752
rect 8236 70688 8252 70752
rect 8316 70688 8324 70752
rect 8004 69664 8324 70688
rect 8004 69600 8012 69664
rect 8076 69600 8092 69664
rect 8156 69600 8172 69664
rect 8236 69600 8252 69664
rect 8316 69600 8324 69664
rect 8004 69354 8324 69600
rect 8004 69118 8046 69354
rect 8282 69118 8324 69354
rect 8004 68576 8324 69118
rect 8004 68512 8012 68576
rect 8076 68512 8092 68576
rect 8156 68512 8172 68576
rect 8236 68512 8252 68576
rect 8316 68512 8324 68576
rect 8004 67488 8324 68512
rect 8004 67424 8012 67488
rect 8076 67424 8092 67488
rect 8156 67424 8172 67488
rect 8236 67424 8252 67488
rect 8316 67424 8324 67488
rect 8004 66400 8324 67424
rect 8004 66336 8012 66400
rect 8076 66336 8092 66400
rect 8156 66336 8172 66400
rect 8236 66336 8252 66400
rect 8316 66336 8324 66400
rect 8004 65312 8324 66336
rect 8004 65248 8012 65312
rect 8076 65248 8092 65312
rect 8156 65248 8172 65312
rect 8236 65248 8252 65312
rect 8316 65248 8324 65312
rect 8004 64354 8324 65248
rect 8004 64224 8046 64354
rect 8282 64224 8324 64354
rect 8004 64160 8012 64224
rect 8316 64160 8324 64224
rect 8004 64118 8046 64160
rect 8282 64118 8324 64160
rect 8004 63136 8324 64118
rect 8004 63072 8012 63136
rect 8076 63072 8092 63136
rect 8156 63072 8172 63136
rect 8236 63072 8252 63136
rect 8316 63072 8324 63136
rect 8004 62048 8324 63072
rect 8004 61984 8012 62048
rect 8076 61984 8092 62048
rect 8156 61984 8172 62048
rect 8236 61984 8252 62048
rect 8316 61984 8324 62048
rect 8004 60960 8324 61984
rect 8004 60896 8012 60960
rect 8076 60896 8092 60960
rect 8156 60896 8172 60960
rect 8236 60896 8252 60960
rect 8316 60896 8324 60960
rect 8004 59872 8324 60896
rect 8004 59808 8012 59872
rect 8076 59808 8092 59872
rect 8156 59808 8172 59872
rect 8236 59808 8252 59872
rect 8316 59808 8324 59872
rect 8004 59354 8324 59808
rect 8004 59118 8046 59354
rect 8282 59118 8324 59354
rect 8004 58784 8324 59118
rect 8004 58720 8012 58784
rect 8076 58720 8092 58784
rect 8156 58720 8172 58784
rect 8236 58720 8252 58784
rect 8316 58720 8324 58784
rect 8004 57696 8324 58720
rect 8004 57632 8012 57696
rect 8076 57632 8092 57696
rect 8156 57632 8172 57696
rect 8236 57632 8252 57696
rect 8316 57632 8324 57696
rect 8004 56608 8324 57632
rect 8004 56544 8012 56608
rect 8076 56544 8092 56608
rect 8156 56544 8172 56608
rect 8236 56544 8252 56608
rect 8316 56544 8324 56608
rect 8004 55520 8324 56544
rect 8004 55456 8012 55520
rect 8076 55456 8092 55520
rect 8156 55456 8172 55520
rect 8236 55456 8252 55520
rect 8316 55456 8324 55520
rect 8004 54432 8324 55456
rect 8004 54368 8012 54432
rect 8076 54368 8092 54432
rect 8156 54368 8172 54432
rect 8236 54368 8252 54432
rect 8316 54368 8324 54432
rect 8004 54354 8324 54368
rect 8004 54118 8046 54354
rect 8282 54118 8324 54354
rect 8004 53344 8324 54118
rect 8004 53280 8012 53344
rect 8076 53280 8092 53344
rect 8156 53280 8172 53344
rect 8236 53280 8252 53344
rect 8316 53280 8324 53344
rect 8004 52256 8324 53280
rect 8004 52192 8012 52256
rect 8076 52192 8092 52256
rect 8156 52192 8172 52256
rect 8236 52192 8252 52256
rect 8316 52192 8324 52256
rect 8004 51168 8324 52192
rect 8004 51104 8012 51168
rect 8076 51104 8092 51168
rect 8156 51104 8172 51168
rect 8236 51104 8252 51168
rect 8316 51104 8324 51168
rect 8004 50080 8324 51104
rect 8004 50016 8012 50080
rect 8076 50016 8092 50080
rect 8156 50016 8172 50080
rect 8236 50016 8252 50080
rect 8316 50016 8324 50080
rect 8004 49354 8324 50016
rect 8004 49118 8046 49354
rect 8282 49118 8324 49354
rect 8004 48992 8324 49118
rect 8004 48928 8012 48992
rect 8076 48928 8092 48992
rect 8156 48928 8172 48992
rect 8236 48928 8252 48992
rect 8316 48928 8324 48992
rect 8004 47904 8324 48928
rect 8004 47840 8012 47904
rect 8076 47840 8092 47904
rect 8156 47840 8172 47904
rect 8236 47840 8252 47904
rect 8316 47840 8324 47904
rect 8004 46816 8324 47840
rect 8004 46752 8012 46816
rect 8076 46752 8092 46816
rect 8156 46752 8172 46816
rect 8236 46752 8252 46816
rect 8316 46752 8324 46816
rect 8004 45728 8324 46752
rect 8004 45664 8012 45728
rect 8076 45664 8092 45728
rect 8156 45664 8172 45728
rect 8236 45664 8252 45728
rect 8316 45664 8324 45728
rect 8004 44640 8324 45664
rect 8004 44576 8012 44640
rect 8076 44576 8092 44640
rect 8156 44576 8172 44640
rect 8236 44576 8252 44640
rect 8316 44576 8324 44640
rect 8004 44354 8324 44576
rect 8004 44118 8046 44354
rect 8282 44118 8324 44354
rect 8004 43552 8324 44118
rect 8004 43488 8012 43552
rect 8076 43488 8092 43552
rect 8156 43488 8172 43552
rect 8236 43488 8252 43552
rect 8316 43488 8324 43552
rect 8004 42464 8324 43488
rect 8004 42400 8012 42464
rect 8076 42400 8092 42464
rect 8156 42400 8172 42464
rect 8236 42400 8252 42464
rect 8316 42400 8324 42464
rect 8004 41376 8324 42400
rect 8004 41312 8012 41376
rect 8076 41312 8092 41376
rect 8156 41312 8172 41376
rect 8236 41312 8252 41376
rect 8316 41312 8324 41376
rect 8004 40288 8324 41312
rect 8004 40224 8012 40288
rect 8076 40224 8092 40288
rect 8156 40224 8172 40288
rect 8236 40224 8252 40288
rect 8316 40224 8324 40288
rect 8004 39354 8324 40224
rect 8004 39200 8046 39354
rect 8282 39200 8324 39354
rect 8004 39136 8012 39200
rect 8316 39136 8324 39200
rect 8004 39118 8046 39136
rect 8282 39118 8324 39136
rect 8004 38112 8324 39118
rect 8004 38048 8012 38112
rect 8076 38048 8092 38112
rect 8156 38048 8172 38112
rect 8236 38048 8252 38112
rect 8316 38048 8324 38112
rect 8004 37024 8324 38048
rect 8004 36960 8012 37024
rect 8076 36960 8092 37024
rect 8156 36960 8172 37024
rect 8236 36960 8252 37024
rect 8316 36960 8324 37024
rect 8004 35936 8324 36960
rect 8004 35872 8012 35936
rect 8076 35872 8092 35936
rect 8156 35872 8172 35936
rect 8236 35872 8252 35936
rect 8316 35872 8324 35936
rect 8004 34848 8324 35872
rect 8004 34784 8012 34848
rect 8076 34784 8092 34848
rect 8156 34784 8172 34848
rect 8236 34784 8252 34848
rect 8316 34784 8324 34848
rect 8004 34354 8324 34784
rect 8004 34118 8046 34354
rect 8282 34118 8324 34354
rect 8004 33760 8324 34118
rect 8004 33696 8012 33760
rect 8076 33696 8092 33760
rect 8156 33696 8172 33760
rect 8236 33696 8252 33760
rect 8316 33696 8324 33760
rect 8004 32672 8324 33696
rect 8004 32608 8012 32672
rect 8076 32608 8092 32672
rect 8156 32608 8172 32672
rect 8236 32608 8252 32672
rect 8316 32608 8324 32672
rect 8004 31584 8324 32608
rect 8004 31520 8012 31584
rect 8076 31520 8092 31584
rect 8156 31520 8172 31584
rect 8236 31520 8252 31584
rect 8316 31520 8324 31584
rect 8004 30496 8324 31520
rect 8004 30432 8012 30496
rect 8076 30432 8092 30496
rect 8156 30432 8172 30496
rect 8236 30432 8252 30496
rect 8316 30432 8324 30496
rect 8004 29408 8324 30432
rect 8004 29344 8012 29408
rect 8076 29354 8092 29408
rect 8156 29354 8172 29408
rect 8236 29354 8252 29408
rect 8316 29344 8324 29408
rect 8004 29118 8046 29344
rect 8282 29118 8324 29344
rect 8004 28320 8324 29118
rect 8004 28256 8012 28320
rect 8076 28256 8092 28320
rect 8156 28256 8172 28320
rect 8236 28256 8252 28320
rect 8316 28256 8324 28320
rect 8004 27232 8324 28256
rect 8004 27168 8012 27232
rect 8076 27168 8092 27232
rect 8156 27168 8172 27232
rect 8236 27168 8252 27232
rect 8316 27168 8324 27232
rect 8004 26144 8324 27168
rect 8004 26080 8012 26144
rect 8076 26080 8092 26144
rect 8156 26080 8172 26144
rect 8236 26080 8252 26144
rect 8316 26080 8324 26144
rect 8004 25056 8324 26080
rect 8004 24992 8012 25056
rect 8076 24992 8092 25056
rect 8156 24992 8172 25056
rect 8236 24992 8252 25056
rect 8316 24992 8324 25056
rect 8004 24354 8324 24992
rect 8004 24118 8046 24354
rect 8282 24118 8324 24354
rect 8004 23968 8324 24118
rect 8004 23904 8012 23968
rect 8076 23904 8092 23968
rect 8156 23904 8172 23968
rect 8236 23904 8252 23968
rect 8316 23904 8324 23968
rect 8004 22880 8324 23904
rect 8004 22816 8012 22880
rect 8076 22816 8092 22880
rect 8156 22816 8172 22880
rect 8236 22816 8252 22880
rect 8316 22816 8324 22880
rect 8004 21792 8324 22816
rect 8004 21728 8012 21792
rect 8076 21728 8092 21792
rect 8156 21728 8172 21792
rect 8236 21728 8252 21792
rect 8316 21728 8324 21792
rect 8004 20704 8324 21728
rect 8004 20640 8012 20704
rect 8076 20640 8092 20704
rect 8156 20640 8172 20704
rect 8236 20640 8252 20704
rect 8316 20640 8324 20704
rect 8004 19616 8324 20640
rect 8004 19552 8012 19616
rect 8076 19552 8092 19616
rect 8156 19552 8172 19616
rect 8236 19552 8252 19616
rect 8316 19552 8324 19616
rect 8004 19354 8324 19552
rect 8004 19118 8046 19354
rect 8282 19118 8324 19354
rect 8004 18528 8324 19118
rect 8004 18464 8012 18528
rect 8076 18464 8092 18528
rect 8156 18464 8172 18528
rect 8236 18464 8252 18528
rect 8316 18464 8324 18528
rect 8004 17440 8324 18464
rect 8004 17376 8012 17440
rect 8076 17376 8092 17440
rect 8156 17376 8172 17440
rect 8236 17376 8252 17440
rect 8316 17376 8324 17440
rect 8004 16352 8324 17376
rect 8004 16288 8012 16352
rect 8076 16288 8092 16352
rect 8156 16288 8172 16352
rect 8236 16288 8252 16352
rect 8316 16288 8324 16352
rect 8004 15264 8324 16288
rect 8004 15200 8012 15264
rect 8076 15200 8092 15264
rect 8156 15200 8172 15264
rect 8236 15200 8252 15264
rect 8316 15200 8324 15264
rect 8004 14354 8324 15200
rect 8004 14176 8046 14354
rect 8282 14176 8324 14354
rect 8004 14112 8012 14176
rect 8076 14112 8092 14118
rect 8156 14112 8172 14118
rect 8236 14112 8252 14118
rect 8316 14112 8324 14176
rect 8004 13088 8324 14112
rect 8004 13024 8012 13088
rect 8076 13024 8092 13088
rect 8156 13024 8172 13088
rect 8236 13024 8252 13088
rect 8316 13024 8324 13088
rect 8004 12000 8324 13024
rect 8004 11936 8012 12000
rect 8076 11936 8092 12000
rect 8156 11936 8172 12000
rect 8236 11936 8252 12000
rect 8316 11936 8324 12000
rect 8004 10912 8324 11936
rect 8004 10848 8012 10912
rect 8076 10848 8092 10912
rect 8156 10848 8172 10912
rect 8236 10848 8252 10912
rect 8316 10848 8324 10912
rect 8004 9824 8324 10848
rect 8004 9760 8012 9824
rect 8076 9760 8092 9824
rect 8156 9760 8172 9824
rect 8236 9760 8252 9824
rect 8316 9760 8324 9824
rect 8004 9354 8324 9760
rect 8004 9118 8046 9354
rect 8282 9118 8324 9354
rect 8004 8736 8324 9118
rect 8004 8672 8012 8736
rect 8076 8672 8092 8736
rect 8156 8672 8172 8736
rect 8236 8672 8252 8736
rect 8316 8672 8324 8736
rect 8004 7648 8324 8672
rect 8004 7584 8012 7648
rect 8076 7584 8092 7648
rect 8156 7584 8172 7648
rect 8236 7584 8252 7648
rect 8316 7584 8324 7648
rect 8004 6560 8324 7584
rect 8004 6496 8012 6560
rect 8076 6496 8092 6560
rect 8156 6496 8172 6560
rect 8236 6496 8252 6560
rect 8316 6496 8324 6560
rect 8004 5472 8324 6496
rect 8004 5408 8012 5472
rect 8076 5408 8092 5472
rect 8156 5408 8172 5472
rect 8236 5408 8252 5472
rect 8316 5408 8324 5472
rect 8004 4384 8324 5408
rect 8004 4320 8012 4384
rect 8076 4354 8092 4384
rect 8156 4354 8172 4384
rect 8236 4354 8252 4384
rect 8316 4320 8324 4384
rect 8004 4118 8046 4320
rect 8282 4118 8324 4320
rect 8004 3296 8324 4118
rect 8004 3232 8012 3296
rect 8076 3232 8092 3296
rect 8156 3232 8172 3296
rect 8236 3232 8252 3296
rect 8316 3232 8324 3296
rect 8004 2208 8324 3232
rect 8004 2144 8012 2208
rect 8076 2144 8092 2208
rect 8156 2144 8172 2208
rect 8236 2144 8252 2208
rect 8316 2144 8324 2208
rect 8004 274 8324 2144
rect 10032 79270 10352 79312
rect 10032 79034 10074 79270
rect 10310 79034 10352 79270
rect 10032 73694 10352 79034
rect 10032 73458 10074 73694
rect 10310 73458 10352 73694
rect 10032 68694 10352 73458
rect 10032 68458 10074 68694
rect 10310 68458 10352 68694
rect 10032 63694 10352 68458
rect 10032 63458 10074 63694
rect 10310 63458 10352 63694
rect 10032 58694 10352 63458
rect 10032 58458 10074 58694
rect 10310 58458 10352 58694
rect 10032 53694 10352 58458
rect 10032 53458 10074 53694
rect 10310 53458 10352 53694
rect 10032 48694 10352 53458
rect 10032 48458 10074 48694
rect 10310 48458 10352 48694
rect 10032 43694 10352 48458
rect 10032 43458 10074 43694
rect 10310 43458 10352 43694
rect 10032 38694 10352 43458
rect 10032 38458 10074 38694
rect 10310 38458 10352 38694
rect 10032 33694 10352 38458
rect 10032 33458 10074 33694
rect 10310 33458 10352 33694
rect 10032 28694 10352 33458
rect 10032 28458 10074 28694
rect 10310 28458 10352 28694
rect 10032 23694 10352 28458
rect 10032 23458 10074 23694
rect 10310 23458 10352 23694
rect 10032 18694 10352 23458
rect 10032 18458 10074 18694
rect 10310 18458 10352 18694
rect 10032 13694 10352 18458
rect 10032 13458 10074 13694
rect 10310 13458 10352 13694
rect 10032 8694 10352 13458
rect 10032 8458 10074 8694
rect 10310 8458 10352 8694
rect 10032 3694 10352 8458
rect 10032 3458 10074 3694
rect 10310 3458 10352 3694
rect 10032 934 10352 3458
rect 10032 698 10074 934
rect 10310 698 10352 934
rect 10032 656 10352 698
rect 10692 74354 11012 79694
rect 10692 74118 10734 74354
rect 10970 74118 11012 74354
rect 10692 69354 11012 74118
rect 10692 69118 10734 69354
rect 10970 69118 11012 69354
rect 10692 64354 11012 69118
rect 10692 64118 10734 64354
rect 10970 64118 11012 64354
rect 10692 59354 11012 64118
rect 10692 59118 10734 59354
rect 10970 59118 11012 59354
rect 10692 54354 11012 59118
rect 10692 54118 10734 54354
rect 10970 54118 11012 54354
rect 10692 49354 11012 54118
rect 10692 49118 10734 49354
rect 10970 49118 11012 49354
rect 10692 44354 11012 49118
rect 10692 44118 10734 44354
rect 10970 44118 11012 44354
rect 10692 39354 11012 44118
rect 10692 39118 10734 39354
rect 10970 39118 11012 39354
rect 10692 34354 11012 39118
rect 10692 34118 10734 34354
rect 10970 34118 11012 34354
rect 10692 29354 11012 34118
rect 10692 29118 10734 29354
rect 10970 29118 11012 29354
rect 10692 24354 11012 29118
rect 10692 24118 10734 24354
rect 10970 24118 11012 24354
rect 10692 19354 11012 24118
rect 10692 19118 10734 19354
rect 10970 19118 11012 19354
rect 10692 14354 11012 19118
rect 10692 14118 10734 14354
rect 10970 14118 11012 14354
rect 10692 9354 11012 14118
rect 10692 9118 10734 9354
rect 10970 9118 11012 9354
rect 10692 4354 11012 9118
rect 10692 4118 10734 4354
rect 10970 4118 11012 4354
rect 8004 38 8046 274
rect 8282 38 8324 274
rect 8004 -4 8324 38
rect 10692 274 11012 4118
rect 10692 38 10734 274
rect 10970 38 11012 274
rect 10692 -4 11012 38
<< via4 >>
rect -1034 79694 -798 79930
rect -1034 74118 -798 74354
rect -1034 69118 -798 69354
rect -1034 64118 -798 64354
rect -1034 59118 -798 59354
rect -1034 54118 -798 54354
rect -1034 49118 -798 49354
rect -1034 44118 -798 44354
rect -1034 39118 -798 39354
rect -1034 34118 -798 34354
rect -1034 29118 -798 29354
rect -1034 24118 -798 24354
rect -1034 19118 -798 19354
rect -1034 14118 -798 14354
rect -1034 9118 -798 9354
rect -1034 4118 -798 4354
rect -374 79034 -138 79270
rect -374 73458 -138 73694
rect -374 68458 -138 68694
rect -374 63458 -138 63694
rect -374 58458 -138 58694
rect -374 53458 -138 53694
rect -374 48458 -138 48694
rect -374 43458 -138 43694
rect -374 38458 -138 38694
rect -374 33458 -138 33694
rect -374 28458 -138 28694
rect -374 23458 -138 23694
rect -374 18458 -138 18694
rect -374 13458 -138 13694
rect -374 8458 -138 8694
rect -374 3458 -138 3694
rect -374 698 -138 934
rect 2386 79034 2622 79270
rect 2386 73472 2622 73694
rect 2386 73458 2416 73472
rect 2416 73458 2432 73472
rect 2432 73458 2496 73472
rect 2496 73458 2512 73472
rect 2512 73458 2576 73472
rect 2576 73458 2592 73472
rect 2592 73458 2622 73472
rect 2386 68458 2622 68694
rect 2386 63680 2622 63694
rect 2386 63616 2416 63680
rect 2416 63616 2432 63680
rect 2432 63616 2496 63680
rect 2496 63616 2512 63680
rect 2512 63616 2576 63680
rect 2576 63616 2592 63680
rect 2592 63616 2622 63680
rect 2386 63458 2622 63616
rect 2386 58458 2622 58694
rect 2386 53458 2622 53694
rect 2386 48458 2622 48694
rect 2386 43458 2622 43694
rect 2386 38656 2622 38694
rect 2386 38592 2416 38656
rect 2416 38592 2432 38656
rect 2432 38592 2496 38656
rect 2496 38592 2512 38656
rect 2512 38592 2576 38656
rect 2576 38592 2592 38656
rect 2592 38592 2622 38656
rect 2386 38458 2622 38592
rect 2386 33458 2622 33694
rect 2386 28458 2622 28694
rect 2386 23458 2622 23694
rect 2386 18458 2622 18694
rect 2386 13632 2622 13694
rect 2386 13568 2416 13632
rect 2416 13568 2432 13632
rect 2432 13568 2496 13632
rect 2496 13568 2512 13632
rect 2512 13568 2576 13632
rect 2576 13568 2592 13632
rect 2592 13568 2622 13632
rect 2386 13458 2622 13568
rect 2386 8458 2622 8694
rect 2386 3458 2622 3694
rect 2386 698 2622 934
rect -1034 38 -798 274
rect 3046 79694 3282 79930
rect 3046 74118 3282 74354
rect 3046 69118 3282 69354
rect 3046 64224 3282 64354
rect 3046 64160 3076 64224
rect 3076 64160 3092 64224
rect 3092 64160 3156 64224
rect 3156 64160 3172 64224
rect 3172 64160 3236 64224
rect 3236 64160 3252 64224
rect 3252 64160 3282 64224
rect 3046 64118 3282 64160
rect 3046 59118 3282 59354
rect 3046 54118 3282 54354
rect 3046 49118 3282 49354
rect 3046 44118 3282 44354
rect 7386 79034 7622 79270
rect 7386 73472 7622 73694
rect 7386 73458 7416 73472
rect 7416 73458 7432 73472
rect 7432 73458 7496 73472
rect 7496 73458 7512 73472
rect 7512 73458 7576 73472
rect 7576 73458 7592 73472
rect 7592 73458 7622 73472
rect 7386 68458 7622 68694
rect 7386 63680 7622 63694
rect 7386 63616 7416 63680
rect 7416 63616 7432 63680
rect 7432 63616 7496 63680
rect 7496 63616 7512 63680
rect 7512 63616 7576 63680
rect 7576 63616 7592 63680
rect 7592 63616 7622 63680
rect 7386 63458 7622 63616
rect 7386 58458 7622 58694
rect 7386 53458 7622 53694
rect 7386 48458 7622 48694
rect 7386 43458 7622 43694
rect 3046 39200 3282 39354
rect 3046 39136 3076 39200
rect 3076 39136 3092 39200
rect 3092 39136 3156 39200
rect 3156 39136 3172 39200
rect 3172 39136 3236 39200
rect 3236 39136 3252 39200
rect 3252 39136 3282 39200
rect 3046 39118 3282 39136
rect 3046 34118 3282 34354
rect 3046 29344 3076 29354
rect 3076 29344 3092 29354
rect 3092 29344 3156 29354
rect 3156 29344 3172 29354
rect 3172 29344 3236 29354
rect 3236 29344 3252 29354
rect 3252 29344 3282 29354
rect 3046 29118 3282 29344
rect 3046 24118 3282 24354
rect 3046 19118 3282 19354
rect 3046 14176 3282 14354
rect 3046 14118 3076 14176
rect 3076 14118 3092 14176
rect 3092 14118 3156 14176
rect 3156 14118 3172 14176
rect 3172 14118 3236 14176
rect 3236 14118 3252 14176
rect 3252 14118 3282 14176
rect 3046 9118 3282 9354
rect 3046 4320 3076 4354
rect 3076 4320 3092 4354
rect 3092 4320 3156 4354
rect 3156 4320 3172 4354
rect 3172 4320 3236 4354
rect 3236 4320 3252 4354
rect 3252 4320 3282 4354
rect 3046 4118 3282 4320
rect 7386 38656 7622 38694
rect 7386 38592 7416 38656
rect 7416 38592 7432 38656
rect 7432 38592 7496 38656
rect 7496 38592 7512 38656
rect 7512 38592 7576 38656
rect 7576 38592 7592 38656
rect 7592 38592 7622 38656
rect 7386 38458 7622 38592
rect 7386 33458 7622 33694
rect 7386 28458 7622 28694
rect 7386 23458 7622 23694
rect 7386 18458 7622 18694
rect 7386 13632 7622 13694
rect 7386 13568 7416 13632
rect 7416 13568 7432 13632
rect 7432 13568 7496 13632
rect 7496 13568 7512 13632
rect 7512 13568 7576 13632
rect 7576 13568 7592 13632
rect 7592 13568 7622 13632
rect 7386 13458 7622 13568
rect 7386 8458 7622 8694
rect 7386 3458 7622 3694
rect 3046 38 3282 274
rect 7386 698 7622 934
rect 8046 79694 8282 79930
rect 10734 79694 10970 79930
rect 8046 74118 8282 74354
rect 8046 69118 8282 69354
rect 8046 64224 8282 64354
rect 8046 64160 8076 64224
rect 8076 64160 8092 64224
rect 8092 64160 8156 64224
rect 8156 64160 8172 64224
rect 8172 64160 8236 64224
rect 8236 64160 8252 64224
rect 8252 64160 8282 64224
rect 8046 64118 8282 64160
rect 8046 59118 8282 59354
rect 8046 54118 8282 54354
rect 8046 49118 8282 49354
rect 8046 44118 8282 44354
rect 8046 39200 8282 39354
rect 8046 39136 8076 39200
rect 8076 39136 8092 39200
rect 8092 39136 8156 39200
rect 8156 39136 8172 39200
rect 8172 39136 8236 39200
rect 8236 39136 8252 39200
rect 8252 39136 8282 39200
rect 8046 39118 8282 39136
rect 8046 34118 8282 34354
rect 8046 29344 8076 29354
rect 8076 29344 8092 29354
rect 8092 29344 8156 29354
rect 8156 29344 8172 29354
rect 8172 29344 8236 29354
rect 8236 29344 8252 29354
rect 8252 29344 8282 29354
rect 8046 29118 8282 29344
rect 8046 24118 8282 24354
rect 8046 19118 8282 19354
rect 8046 14176 8282 14354
rect 8046 14118 8076 14176
rect 8076 14118 8092 14176
rect 8092 14118 8156 14176
rect 8156 14118 8172 14176
rect 8172 14118 8236 14176
rect 8236 14118 8252 14176
rect 8252 14118 8282 14176
rect 8046 9118 8282 9354
rect 8046 4320 8076 4354
rect 8076 4320 8092 4354
rect 8092 4320 8156 4354
rect 8156 4320 8172 4354
rect 8172 4320 8236 4354
rect 8236 4320 8252 4354
rect 8252 4320 8282 4354
rect 8046 4118 8282 4320
rect 10074 79034 10310 79270
rect 10074 73458 10310 73694
rect 10074 68458 10310 68694
rect 10074 63458 10310 63694
rect 10074 58458 10310 58694
rect 10074 53458 10310 53694
rect 10074 48458 10310 48694
rect 10074 43458 10310 43694
rect 10074 38458 10310 38694
rect 10074 33458 10310 33694
rect 10074 28458 10310 28694
rect 10074 23458 10310 23694
rect 10074 18458 10310 18694
rect 10074 13458 10310 13694
rect 10074 8458 10310 8694
rect 10074 3458 10310 3694
rect 10074 698 10310 934
rect 10734 74118 10970 74354
rect 10734 69118 10970 69354
rect 10734 64118 10970 64354
rect 10734 59118 10970 59354
rect 10734 54118 10970 54354
rect 10734 49118 10970 49354
rect 10734 44118 10970 44354
rect 10734 39118 10970 39354
rect 10734 34118 10970 34354
rect 10734 29118 10970 29354
rect 10734 24118 10970 24354
rect 10734 19118 10970 19354
rect 10734 14118 10970 14354
rect 10734 9118 10970 9354
rect 10734 4118 10970 4354
rect 8046 38 8282 274
rect 10734 38 10970 274
<< metal5 >>
rect -1076 79930 11012 79972
rect -1076 79694 -1034 79930
rect -798 79694 3046 79930
rect 3282 79694 8046 79930
rect 8282 79694 10734 79930
rect 10970 79694 11012 79930
rect -1076 79652 11012 79694
rect -416 79270 10352 79312
rect -416 79034 -374 79270
rect -138 79034 2386 79270
rect 2622 79034 7386 79270
rect 7622 79034 10074 79270
rect 10310 79034 10352 79270
rect -416 78992 10352 79034
rect -1076 74354 11012 74396
rect -1076 74118 -1034 74354
rect -798 74118 3046 74354
rect 3282 74118 8046 74354
rect 8282 74118 10734 74354
rect 10970 74118 11012 74354
rect -1076 74076 11012 74118
rect -1076 73694 11012 73736
rect -1076 73458 -374 73694
rect -138 73458 2386 73694
rect 2622 73458 7386 73694
rect 7622 73458 10074 73694
rect 10310 73458 11012 73694
rect -1076 73416 11012 73458
rect -1076 69354 11012 69396
rect -1076 69118 -1034 69354
rect -798 69118 3046 69354
rect 3282 69118 8046 69354
rect 8282 69118 10734 69354
rect 10970 69118 11012 69354
rect -1076 69076 11012 69118
rect -1076 68694 11012 68736
rect -1076 68458 -374 68694
rect -138 68458 2386 68694
rect 2622 68458 7386 68694
rect 7622 68458 10074 68694
rect 10310 68458 11012 68694
rect -1076 68416 11012 68458
rect -1076 64354 11012 64396
rect -1076 64118 -1034 64354
rect -798 64118 3046 64354
rect 3282 64118 8046 64354
rect 8282 64118 10734 64354
rect 10970 64118 11012 64354
rect -1076 64076 11012 64118
rect -1076 63694 11012 63736
rect -1076 63458 -374 63694
rect -138 63458 2386 63694
rect 2622 63458 7386 63694
rect 7622 63458 10074 63694
rect 10310 63458 11012 63694
rect -1076 63416 11012 63458
rect -1076 59354 11012 59396
rect -1076 59118 -1034 59354
rect -798 59118 3046 59354
rect 3282 59118 8046 59354
rect 8282 59118 10734 59354
rect 10970 59118 11012 59354
rect -1076 59076 11012 59118
rect -1076 58694 11012 58736
rect -1076 58458 -374 58694
rect -138 58458 2386 58694
rect 2622 58458 7386 58694
rect 7622 58458 10074 58694
rect 10310 58458 11012 58694
rect -1076 58416 11012 58458
rect -1076 54354 11012 54396
rect -1076 54118 -1034 54354
rect -798 54118 3046 54354
rect 3282 54118 8046 54354
rect 8282 54118 10734 54354
rect 10970 54118 11012 54354
rect -1076 54076 11012 54118
rect -1076 53694 11012 53736
rect -1076 53458 -374 53694
rect -138 53458 2386 53694
rect 2622 53458 7386 53694
rect 7622 53458 10074 53694
rect 10310 53458 11012 53694
rect -1076 53416 11012 53458
rect -1076 49354 11012 49396
rect -1076 49118 -1034 49354
rect -798 49118 3046 49354
rect 3282 49118 8046 49354
rect 8282 49118 10734 49354
rect 10970 49118 11012 49354
rect -1076 49076 11012 49118
rect -1076 48694 11012 48736
rect -1076 48458 -374 48694
rect -138 48458 2386 48694
rect 2622 48458 7386 48694
rect 7622 48458 10074 48694
rect 10310 48458 11012 48694
rect -1076 48416 11012 48458
rect -1076 44354 11012 44396
rect -1076 44118 -1034 44354
rect -798 44118 3046 44354
rect 3282 44118 8046 44354
rect 8282 44118 10734 44354
rect 10970 44118 11012 44354
rect -1076 44076 11012 44118
rect -1076 43694 11012 43736
rect -1076 43458 -374 43694
rect -138 43458 2386 43694
rect 2622 43458 7386 43694
rect 7622 43458 10074 43694
rect 10310 43458 11012 43694
rect -1076 43416 11012 43458
rect -1076 39354 11012 39396
rect -1076 39118 -1034 39354
rect -798 39118 3046 39354
rect 3282 39118 8046 39354
rect 8282 39118 10734 39354
rect 10970 39118 11012 39354
rect -1076 39076 11012 39118
rect -1076 38694 11012 38736
rect -1076 38458 -374 38694
rect -138 38458 2386 38694
rect 2622 38458 7386 38694
rect 7622 38458 10074 38694
rect 10310 38458 11012 38694
rect -1076 38416 11012 38458
rect -1076 34354 11012 34396
rect -1076 34118 -1034 34354
rect -798 34118 3046 34354
rect 3282 34118 8046 34354
rect 8282 34118 10734 34354
rect 10970 34118 11012 34354
rect -1076 34076 11012 34118
rect -1076 33694 11012 33736
rect -1076 33458 -374 33694
rect -138 33458 2386 33694
rect 2622 33458 7386 33694
rect 7622 33458 10074 33694
rect 10310 33458 11012 33694
rect -1076 33416 11012 33458
rect -1076 29354 11012 29396
rect -1076 29118 -1034 29354
rect -798 29118 3046 29354
rect 3282 29118 8046 29354
rect 8282 29118 10734 29354
rect 10970 29118 11012 29354
rect -1076 29076 11012 29118
rect -1076 28694 11012 28736
rect -1076 28458 -374 28694
rect -138 28458 2386 28694
rect 2622 28458 7386 28694
rect 7622 28458 10074 28694
rect 10310 28458 11012 28694
rect -1076 28416 11012 28458
rect -1076 24354 11012 24396
rect -1076 24118 -1034 24354
rect -798 24118 3046 24354
rect 3282 24118 8046 24354
rect 8282 24118 10734 24354
rect 10970 24118 11012 24354
rect -1076 24076 11012 24118
rect -1076 23694 11012 23736
rect -1076 23458 -374 23694
rect -138 23458 2386 23694
rect 2622 23458 7386 23694
rect 7622 23458 10074 23694
rect 10310 23458 11012 23694
rect -1076 23416 11012 23458
rect -1076 19354 11012 19396
rect -1076 19118 -1034 19354
rect -798 19118 3046 19354
rect 3282 19118 8046 19354
rect 8282 19118 10734 19354
rect 10970 19118 11012 19354
rect -1076 19076 11012 19118
rect -1076 18694 11012 18736
rect -1076 18458 -374 18694
rect -138 18458 2386 18694
rect 2622 18458 7386 18694
rect 7622 18458 10074 18694
rect 10310 18458 11012 18694
rect -1076 18416 11012 18458
rect -1076 14354 11012 14396
rect -1076 14118 -1034 14354
rect -798 14118 3046 14354
rect 3282 14118 8046 14354
rect 8282 14118 10734 14354
rect 10970 14118 11012 14354
rect -1076 14076 11012 14118
rect -1076 13694 11012 13736
rect -1076 13458 -374 13694
rect -138 13458 2386 13694
rect 2622 13458 7386 13694
rect 7622 13458 10074 13694
rect 10310 13458 11012 13694
rect -1076 13416 11012 13458
rect -1076 9354 11012 9396
rect -1076 9118 -1034 9354
rect -798 9118 3046 9354
rect 3282 9118 8046 9354
rect 8282 9118 10734 9354
rect 10970 9118 11012 9354
rect -1076 9076 11012 9118
rect -1076 8694 11012 8736
rect -1076 8458 -374 8694
rect -138 8458 2386 8694
rect 2622 8458 7386 8694
rect 7622 8458 10074 8694
rect 10310 8458 11012 8694
rect -1076 8416 11012 8458
rect -1076 4354 11012 4396
rect -1076 4118 -1034 4354
rect -798 4118 3046 4354
rect 3282 4118 8046 4354
rect 8282 4118 10734 4354
rect 10970 4118 11012 4354
rect -1076 4076 11012 4118
rect -1076 3694 11012 3736
rect -1076 3458 -374 3694
rect -138 3458 2386 3694
rect 2622 3458 7386 3694
rect 7622 3458 10074 3694
rect 10310 3458 11012 3694
rect -1076 3416 11012 3458
rect -416 934 10352 976
rect -416 698 -374 934
rect -138 698 2386 934
rect 2622 698 7386 934
rect 7622 698 10074 934
rect 10310 698 10352 934
rect -416 656 10352 698
rect -1076 274 11012 316
rect -1076 38 -1034 274
rect -798 38 3046 274
rect 3282 38 8046 274
rect 8282 38 10734 274
rect 10970 38 11012 274
rect -1076 -4 11012 38
use sky130_fd_sc_hd__mux2_1  _177_
timestamp 1699142937
transform -1 0 8556 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1699142937
transform -1 0 8372 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _179_
timestamp 1699142937
transform -1 0 5152 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1699142937
transform -1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _181_
timestamp 1699142937
transform -1 0 6532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1699142937
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1699142937
transform 1 0 7728 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1699142937
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1699142937
transform 1 0 7728 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1699142937
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1699142937
transform 1 0 7728 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1699142937
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _189_
timestamp 1699142937
transform 1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1699142937
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _191_
timestamp 1699142937
transform 1 0 7728 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1699142937
transform 1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1699142937
transform 1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1699142937
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1699142937
transform 1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1699142937
transform 1 0 6900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _197_
timestamp 1699142937
transform 1 0 7728 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1699142937
transform -1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 1699142937
transform 1 0 7728 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1699142937
transform 1 0 6808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 1699142937
transform 1 0 7728 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1699142937
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 1699142937
transform 1 0 7728 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1699142937
transform 1 0 6808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1699142937
transform 1 0 7728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1699142937
transform 1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1699142937
transform 1 0 7728 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1699142937
transform -1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1699142937
transform 1 0 7728 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1699142937
transform -1 0 6716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1699142937
transform 1 0 7728 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1699142937
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1699142937
transform -1 0 8188 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1699142937
transform 1 0 8188 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _215_
timestamp 1699142937
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1699142937
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _217_
timestamp 1699142937
transform -1 0 6072 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 1699142937
transform 1 0 5244 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _219_
timestamp 1699142937
transform -1 0 7084 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _220_
timestamp 1699142937
transform -1 0 7636 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1699142937
transform 1 0 7544 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1699142937
transform 1 0 6992 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1699142937
transform 1 0 6716 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1699142937
transform -1 0 6716 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1699142937
transform 1 0 6624 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1699142937
transform -1 0 6716 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1699142937
transform 1 0 6716 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1699142937
transform -1 0 6716 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1699142937
transform -1 0 7544 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1699142937
transform 1 0 7544 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1699142937
transform 1 0 6716 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1699142937
transform -1 0 6716 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1699142937
transform -1 0 7636 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1699142937
transform 1 0 7636 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1699142937
transform 1 0 6808 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1699142937
transform -1 0 6716 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1699142937
transform 1 0 6716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1699142937
transform -1 0 6716 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1699142937
transform 1 0 6716 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1699142937
transform -1 0 6716 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _241_
timestamp 1699142937
transform 1 0 7728 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1699142937
transform 1 0 7636 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1699142937
transform -1 0 6716 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1699142937
transform -1 0 7636 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1699142937
transform 1 0 7176 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _246_
timestamp 1699142937
transform 1 0 6808 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1699142937
transform -1 0 6716 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _248_
timestamp 1699142937
transform 1 0 6900 0 1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1699142937
transform 1 0 6992 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _250_
timestamp 1699142937
transform 1 0 7176 0 -1 71808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1699142937
transform 1 0 7176 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _252_
timestamp 1699142937
transform -1 0 7728 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1699142937
transform 1 0 7728 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1699142937
transform 1 0 6900 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1699142937
transform 1 0 6992 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _256_
timestamp 1699142937
transform 1 0 6808 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1699142937
transform -1 0 6716 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1699142937
transform 1 0 6808 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1699142937
transform -1 0 6716 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1699142937
transform -1 0 7636 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1699142937
transform 1 0 7452 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _262_
timestamp 1699142937
transform -1 0 7636 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1699142937
transform 1 0 6624 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1699142937
transform -1 0 6716 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1699142937
transform 1 0 6624 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1699142937
transform -1 0 6716 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1699142937
transform 1 0 6624 0 1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1699142937
transform -1 0 6716 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _269_
timestamp 1699142937
transform 1 0 6624 0 1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1699142937
transform -1 0 6716 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1699142937
transform 1 0 6624 0 -1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1699142937
transform -1 0 6716 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1699142937
transform 1 0 6716 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1699142937
transform -1 0 7084 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1699142937
transform 1 0 6716 0 1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1699142937
transform -1 0 6716 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _277_
timestamp 1699142937
transform 1 0 6716 0 1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1699142937
transform -1 0 6716 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp 1699142937
transform 1 0 6624 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1699142937
transform -1 0 7084 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1699142937
transform 1 0 6716 0 -1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1699142937
transform -1 0 6716 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _283_
timestamp 1699142937
transform 1 0 6348 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1699142937
transform -1 0 6716 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _285_
timestamp 1699142937
transform 1 0 7176 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1699142937
transform -1 0 7084 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1699142937
transform -1 0 7360 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1699142937
transform 1 0 7084 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1699142937
transform 1 0 5428 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1699142937
transform 1 0 5612 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1699142937
transform 1 0 5428 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1699142937
transform 1 0 5060 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1699142937
transform 1 0 5336 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1699142937
transform 1 0 5060 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1699142937
transform 1 0 5428 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1699142937
transform 1 0 5060 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1699142937
transform 1 0 5428 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1699142937
transform 1 0 5152 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1699142937
transform 1 0 5520 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1699142937
transform 1 0 4876 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1699142937
transform 1 0 5428 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1699142937
transform 1 0 5152 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1699142937
transform 1 0 6348 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1699142937
transform 1 0 5152 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _305_
timestamp 1699142937
transform 1 0 5520 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1699142937
transform 1 0 5060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1699142937
transform 1 0 6900 0 1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1699142937
transform 1 0 5612 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1699142937
transform 1 0 6348 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1699142937
transform 1 0 5244 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1699142937
transform 1 0 5428 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1699142937
transform 1 0 5152 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1699142937
transform 1 0 5520 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1699142937
transform 1 0 5152 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1699142937
transform 1 0 5520 0 1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1699142937
transform 1 0 5152 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _317_
timestamp 1699142937
transform 1 0 6348 0 -1 71808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1699142937
transform 1 0 5244 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1699142937
transform 1 0 6348 0 -1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1699142937
transform 1 0 5428 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1699142937
transform 1 0 5520 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1699142937
transform 1 0 5244 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _323_
timestamp 1699142937
transform 1 0 5428 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1699142937
transform 1 0 5152 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp 1699142937
transform 1 0 5428 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1699142937
transform 1 0 5152 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _327_
timestamp 1699142937
transform 1 0 5428 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1699142937
transform 1 0 5060 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1699142937
transform 1 0 5336 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1699142937
transform 1 0 4968 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1699142937
transform 1 0 5244 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1699142937
transform 1 0 4876 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1699142937
transform 1 0 5244 0 1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1699142937
transform 1 0 4968 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1699142937
transform 1 0 5244 0 -1 54400
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1699142937
transform 1 0 4968 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1699142937
transform 1 0 5244 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1699142937
transform 1 0 4968 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1699142937
transform 1 0 5060 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1699142937
transform 1 0 4784 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1699142937
transform 1 0 5244 0 1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1699142937
transform 1 0 4968 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1699142937
transform 1 0 5152 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1699142937
transform 1 0 4876 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1699142937
transform 1 0 5152 0 -1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1699142937
transform 1 0 4784 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1699142937
transform 1 0 5152 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1699142937
transform 1 0 4784 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1699142937
transform 1 0 5244 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1699142937
transform 1 0 4784 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1699142937
transform 1 0 5336 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1699142937
transform 1 0 5152 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1699142937
transform 1 0 5244 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1699142937
transform 1 0 4600 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _355_
timestamp 1699142937
transform 1 0 4692 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 1699142937
transform 1 0 6716 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _357_
timestamp 1699142937
transform 1 0 6716 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _358_
timestamp 1699142937
transform 1 0 6716 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _359_
timestamp 1699142937
transform 1 0 6716 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _360_
timestamp 1699142937
transform 1 0 6716 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _361_
timestamp 1699142937
transform 1 0 6716 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _362_
timestamp 1699142937
transform 1 0 6716 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _363_
timestamp 1699142937
transform 1 0 6716 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 1699142937
transform 1 0 6716 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _365_
timestamp 1699142937
transform 1 0 6716 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp 1699142937
transform 1 0 6716 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp 1699142937
transform 1 0 6716 0 1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp 1699142937
transform 1 0 6716 0 1 68544
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _369_
timestamp 1699142937
transform 1 0 6716 0 -1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _370_
timestamp 1699142937
transform 1 0 6716 0 1 71808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp 1699142937
transform 1 0 6716 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _372_
timestamp 1699142937
transform 1 0 6716 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _373_
timestamp 1699142937
transform 1 0 6716 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _374_
timestamp 1699142937
transform 1 0 6716 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _375_
timestamp 1699142937
transform 1 0 6716 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _376_
timestamp 1699142937
transform 1 0 6716 0 1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _377_
timestamp 1699142937
transform 1 0 6716 0 1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _378_
timestamp 1699142937
transform 1 0 6716 0 -1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _379_
timestamp 1699142937
transform 1 0 6716 0 -1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _380_
timestamp 1699142937
transform 1 0 6716 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1699142937
transform 1 0 6716 0 1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1699142937
transform 1 0 6716 0 -1 58752
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1699142937
transform 1 0 6716 0 -1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1699142937
transform 1 0 6716 0 -1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _385_
timestamp 1699142937
transform 1 0 6716 0 1 62016
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _386_
timestamp 1699142937
transform 1 0 6440 0 -1 64192
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _387_
timestamp 1699142937
transform 1 0 6716 0 1 64192
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _388_
timestamp 1699142937
transform 1 0 6532 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1699142937
transform 1 0 3772 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1699142937
transform 1 0 3956 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _391_
timestamp 1699142937
transform 1 0 5152 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _392_
timestamp 1699142937
transform 1 0 6624 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _393_
timestamp 1699142937
transform 1 0 6532 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _394_
timestamp 1699142937
transform 1 0 6532 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _395_
timestamp 1699142937
transform 1 0 6532 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1699142937
transform 1 0 6532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1699142937
transform 1 0 6532 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1699142937
transform -1 0 8372 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1699142937
transform 1 0 6532 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1699142937
transform 1 0 6532 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1699142937
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1699142937
transform 1 0 6532 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1699142937
transform -1 0 8372 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _404_
timestamp 1699142937
transform 1 0 6532 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _405_
timestamp 1699142937
transform 1 0 6532 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _406_
timestamp 1699142937
transform -1 0 8464 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _407_
timestamp 1699142937
transform 1 0 5888 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _408_
timestamp 1699142937
transform 1 0 4048 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _409_
timestamp 1699142937
transform 1 0 4784 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _410_
timestamp 1699142937
transform 1 0 4600 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _411_
timestamp 1699142937
transform 1 0 4416 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _412_
timestamp 1699142937
transform 1 0 4600 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp 1699142937
transform 1 0 4692 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _414_
timestamp 1699142937
transform 1 0 4416 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _415_
timestamp 1699142937
transform 1 0 4784 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _416_
timestamp 1699142937
transform 1 0 4784 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _417_
timestamp 1699142937
transform 1 0 4416 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _418_
timestamp 1699142937
transform 1 0 4784 0 1 65280
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _419_
timestamp 1699142937
transform 1 0 4784 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _420_
timestamp 1699142937
transform 1 0 4784 0 1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _421_
timestamp 1699142937
transform 1 0 4416 0 -1 69632
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _422_
timestamp 1699142937
transform 1 0 4416 0 -1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _423_
timestamp 1699142937
transform 1 0 4784 0 1 71808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1699142937
transform 1 0 5060 0 1 72896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _425_
timestamp 1699142937
transform 1 0 4324 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1699142937
transform 1 0 4416 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1699142937
transform 1 0 4416 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _428_
timestamp 1699142937
transform 1 0 4692 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1699142937
transform 1 0 4508 0 1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _430_
timestamp 1699142937
transform 1 0 4416 0 -1 52224
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _431_
timestamp 1699142937
transform 1 0 4416 0 -1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _432_
timestamp 1699142937
transform 1 0 4508 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1699142937
transform 1 0 4508 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _434_
timestamp 1699142937
transform 1 0 4416 0 -1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1699142937
transform 1 0 4416 0 -1 58752
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _436_
timestamp 1699142937
transform 1 0 4416 0 -1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _437_
timestamp 1699142937
transform 1 0 4416 0 1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _438_
timestamp 1699142937
transform 1 0 4324 0 1 62016
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _439_
timestamp 1699142937
transform 1 0 4324 0 1 63104
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _440_
timestamp 1699142937
transform 1 0 4876 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp 1699142937
transform 1 0 4416 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _442__74
timestamp 1699608013
transform -1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _442_
timestamp 1699142937
transform -1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _443__75
timestamp 1699608013
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _443_
timestamp 1699142937
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1699142937
transform -1 0 5520 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1699142937
transform 1 0 5888 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1699142937
transform -1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1699142937
transform -1 0 6716 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_0_0_clk
timestamp 1699142937
transform 1 0 4600 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_1_0_clk
timestamp 1699142937
transform 1 0 6808 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_2_0_clk
timestamp 1699142937
transform -1 0 6900 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_3_0_clk
timestamp 1699142937
transform 1 0 7268 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_4_0_clk
timestamp 1699142937
transform -1 0 5520 0 -1 50048
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_5_0_clk
timestamp 1699142937
transform -1 0 5612 0 -1 65280
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_6_0_clk
timestamp 1699142937
transform -1 0 7544 0 -1 50048
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_3_7_0_clk
timestamp 1699142937
transform 1 0 6624 0 1 66368
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 1699142937
transform -1 0 7728 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 1699142937
transform 1 0 6716 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1699142937
transform 1 0 7544 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1699142937
transform 1 0 6440 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1699142937
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp 1699142937
transform -1 0 6808 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1699142937
transform 1 0 8004 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1699142937
transform 1 0 6348 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 1699142937
transform 1 0 8004 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 1699142937
transform 1 0 8004 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1699142937
transform 1 0 6348 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1699142937
transform 1 0 7176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 1699142937
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1699142937
transform 1 0 7176 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1699142937
transform -1 0 7820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout71
timestamp 1699142937
transform 1 0 6348 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 1699142937
transform 1 0 6072 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 1699142937
transform -1 0 6348 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_3
timestamp 1699142937
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_9
timestamp 1699142937
transform 1 0 1932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_17
timestamp 1699142937
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 1699142937
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29
timestamp 1699142937
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_38
timestamp 1699142937
transform 1 0 4600 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_46
timestamp 1699142937
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1699142937
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_67
timestamp 1699142937
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1699142937
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1699142937
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_17
timestamp 1699142937
transform 1 0 2668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_25
timestamp 1699142937
transform 1 0 3404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_33
timestamp 1699142937
transform 1 0 4140 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_41
timestamp 1699142937
transform 1 0 4876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_49
timestamp 1699142937
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1699142937
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 1699142937
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_65
timestamp 1699142937
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_73
timestamp 1699142937
transform 1 0 7820 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_3
timestamp 1699142937
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_11
timestamp 1699142937
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1699142937
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1699142937
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1699142937
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_37
timestamp 1699142937
transform 1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_45
timestamp 1699142937
transform 1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1699142937
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_61
timestamp 1699142937
transform 1 0 6716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_69
timestamp 1699142937
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_77
timestamp 1699142937
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1699142937
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_11
timestamp 1699142937
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_19
timestamp 1699142937
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_27
timestamp 1699142937
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_35
timestamp 1699142937
transform 1 0 4324 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_43
timestamp 1699142937
transform 1 0 5060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1699142937
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1699142937
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1699142937
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_65
timestamp 1699142937
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_73
timestamp 1699142937
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 1699142937
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_11
timestamp 1699142937
transform 1 0 2116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1699142937
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1699142937
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1699142937
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_37
timestamp 1699142937
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_45
timestamp 1699142937
transform 1 0 5244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1699142937
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_61
timestamp 1699142937
transform 1 0 6716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_69
timestamp 1699142937
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_77
timestamp 1699142937
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1699142937
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_11
timestamp 1699142937
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_19
timestamp 1699142937
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 1699142937
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_35
timestamp 1699142937
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_43
timestamp 1699142937
transform 1 0 5060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1699142937
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1699142937
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1699142937
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_65
timestamp 1699142937
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_73
timestamp 1699142937
transform 1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1699142937
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_11
timestamp 1699142937
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 1699142937
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1699142937
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1699142937
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_37
timestamp 1699142937
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_45
timestamp 1699142937
transform 1 0 5244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 1699142937
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_61
timestamp 1699142937
transform 1 0 6716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_69
timestamp 1699142937
transform 1 0 7452 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_77
timestamp 1699142937
transform 1 0 8188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1699142937
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_11
timestamp 1699142937
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_19
timestamp 1699142937
transform 1 0 2852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_27
timestamp 1699142937
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_35
timestamp 1699142937
transform 1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_43
timestamp 1699142937
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1699142937
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1699142937
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1699142937
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_65
timestamp 1699142937
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1699142937
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_11
timestamp 1699142937
transform 1 0 2116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_19
timestamp 1699142937
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1699142937
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_49
timestamp 1699142937
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_59
timestamp 1699142937
transform 1 0 6532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_65
timestamp 1699142937
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1699142937
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_11
timestamp 1699142937
transform 1 0 2116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_19
timestamp 1699142937
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1699142937
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_51
timestamp 1699142937
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1699142937
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_80
timestamp 1699142937
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1699142937
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_11
timestamp 1699142937
transform 1 0 2116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 1699142937
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1699142937
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 1699142937
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_35
timestamp 1699142937
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1699142937
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_11
timestamp 1699142937
transform 1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_19
timestamp 1699142937
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_27
timestamp 1699142937
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_35
timestamp 1699142937
transform 1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_43
timestamp 1699142937
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1699142937
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1699142937
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_79
timestamp 1699142937
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1699142937
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_11
timestamp 1699142937
transform 1 0 2116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_19
timestamp 1699142937
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1699142937
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1699142937
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_37
timestamp 1699142937
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_45
timestamp 1699142937
transform 1 0 5244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_53
timestamp 1699142937
transform 1 0 5980 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1699142937
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_11
timestamp 1699142937
transform 1 0 2116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_19
timestamp 1699142937
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_27
timestamp 1699142937
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_35
timestamp 1699142937
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_43
timestamp 1699142937
transform 1 0 5060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1699142937
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1699142937
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1699142937
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_65
timestamp 1699142937
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1699142937
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_11
timestamp 1699142937
transform 1 0 2116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1699142937
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1699142937
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1699142937
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_37
timestamp 1699142937
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_45
timestamp 1699142937
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_53
timestamp 1699142937
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_79
timestamp 1699142937
transform 1 0 8372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1699142937
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_11
timestamp 1699142937
transform 1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_19
timestamp 1699142937
transform 1 0 2852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1699142937
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_35
timestamp 1699142937
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_43
timestamp 1699142937
transform 1 0 5060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1699142937
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1699142937
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1699142937
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1699142937
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_69
timestamp 1699142937
transform 1 0 7452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1699142937
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_11
timestamp 1699142937
transform 1 0 2116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_19
timestamp 1699142937
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1699142937
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1699142937
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_37
timestamp 1699142937
transform 1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_45
timestamp 1699142937
transform 1 0 5244 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_53
timestamp 1699142937
transform 1 0 5980 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_79
timestamp 1699142937
transform 1 0 8372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1699142937
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_11
timestamp 1699142937
transform 1 0 2116 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_19
timestamp 1699142937
transform 1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1699142937
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_35
timestamp 1699142937
transform 1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_43
timestamp 1699142937
transform 1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1699142937
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1699142937
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1699142937
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1699142937
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_11
timestamp 1699142937
transform 1 0 2116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_19
timestamp 1699142937
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1699142937
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1699142937
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_37
timestamp 1699142937
transform 1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_45
timestamp 1699142937
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_53
timestamp 1699142937
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_61
timestamp 1699142937
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1699142937
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_11
timestamp 1699142937
transform 1 0 2116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_19
timestamp 1699142937
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_27
timestamp 1699142937
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_35
timestamp 1699142937
transform 1 0 4324 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_43
timestamp 1699142937
transform 1 0 5060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1699142937
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1699142937
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1699142937
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_79
timestamp 1699142937
transform 1 0 8372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1699142937
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_11
timestamp 1699142937
transform 1 0 2116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 1699142937
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1699142937
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1699142937
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_37
timestamp 1699142937
transform 1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_45
timestamp 1699142937
transform 1 0 5244 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_53
timestamp 1699142937
transform 1 0 5980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1699142937
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1699142937
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_11
timestamp 1699142937
transform 1 0 2116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_19
timestamp 1699142937
transform 1 0 2852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_27
timestamp 1699142937
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_35
timestamp 1699142937
transform 1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_43
timestamp 1699142937
transform 1 0 5060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1699142937
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1699142937
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1699142937
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_79
timestamp 1699142937
transform 1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_3
timestamp 1699142937
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_11
timestamp 1699142937
transform 1 0 2116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_19
timestamp 1699142937
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1699142937
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1699142937
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_37
timestamp 1699142937
transform 1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_45
timestamp 1699142937
transform 1 0 5244 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_51
timestamp 1699142937
transform 1 0 5796 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1699142937
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_11
timestamp 1699142937
transform 1 0 2116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_19
timestamp 1699142937
transform 1 0 2852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_27
timestamp 1699142937
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_35
timestamp 1699142937
transform 1 0 4324 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_43
timestamp 1699142937
transform 1 0 5060 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1699142937
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1699142937
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1699142937
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 1699142937
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_11
timestamp 1699142937
transform 1 0 2116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_19
timestamp 1699142937
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1699142937
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1699142937
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_37
timestamp 1699142937
transform 1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_45
timestamp 1699142937
transform 1 0 5244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_53
timestamp 1699142937
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_79
timestamp 1699142937
transform 1 0 8372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1699142937
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_11
timestamp 1699142937
transform 1 0 2116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_19
timestamp 1699142937
transform 1 0 2852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_27
timestamp 1699142937
transform 1 0 3588 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_35
timestamp 1699142937
transform 1 0 4324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_43
timestamp 1699142937
transform 1 0 5060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1699142937
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1699142937
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_57
timestamp 1699142937
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_65
timestamp 1699142937
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_69
timestamp 1699142937
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1699142937
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_11
timestamp 1699142937
transform 1 0 2116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_19
timestamp 1699142937
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1699142937
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 1699142937
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_37
timestamp 1699142937
transform 1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_45
timestamp 1699142937
transform 1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_53
timestamp 1699142937
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_79
timestamp 1699142937
transform 1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1699142937
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_11
timestamp 1699142937
transform 1 0 2116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_19
timestamp 1699142937
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_27
timestamp 1699142937
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_35
timestamp 1699142937
transform 1 0 4324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_43
timestamp 1699142937
transform 1 0 5060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1699142937
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1699142937
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1699142937
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_3
timestamp 1699142937
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_11
timestamp 1699142937
transform 1 0 2116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_19
timestamp 1699142937
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1699142937
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp 1699142937
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_37
timestamp 1699142937
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_45
timestamp 1699142937
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_53
timestamp 1699142937
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_61
timestamp 1699142937
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1699142937
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_11
timestamp 1699142937
transform 1 0 2116 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_19
timestamp 1699142937
transform 1 0 2852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_27
timestamp 1699142937
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_35
timestamp 1699142937
transform 1 0 4324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_43
timestamp 1699142937
transform 1 0 5060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1699142937
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1699142937
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_57
timestamp 1699142937
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_79
timestamp 1699142937
transform 1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1699142937
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_11
timestamp 1699142937
transform 1 0 2116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_19
timestamp 1699142937
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1699142937
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1699142937
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_37
timestamp 1699142937
transform 1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_45
timestamp 1699142937
transform 1 0 5244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_53
timestamp 1699142937
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_61
timestamp 1699142937
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_65
timestamp 1699142937
transform 1 0 7084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_69
timestamp 1699142937
transform 1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp 1699142937
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_11
timestamp 1699142937
transform 1 0 2116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_19
timestamp 1699142937
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_27
timestamp 1699142937
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_35
timestamp 1699142937
transform 1 0 4324 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_43
timestamp 1699142937
transform 1 0 5060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1699142937
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1699142937
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_57
timestamp 1699142937
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_79
timestamp 1699142937
transform 1 0 8372 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_3
timestamp 1699142937
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_11
timestamp 1699142937
transform 1 0 2116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 1699142937
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1699142937
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1699142937
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_37
timestamp 1699142937
transform 1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_45
timestamp 1699142937
transform 1 0 5244 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_53
timestamp 1699142937
transform 1 0 5980 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1699142937
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_11
timestamp 1699142937
transform 1 0 2116 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_19
timestamp 1699142937
transform 1 0 2852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_27
timestamp 1699142937
transform 1 0 3588 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_35
timestamp 1699142937
transform 1 0 4324 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_43
timestamp 1699142937
transform 1 0 5060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1699142937
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1699142937
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1699142937
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_65
timestamp 1699142937
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 1699142937
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_11
timestamp 1699142937
transform 1 0 2116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1699142937
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1699142937
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1699142937
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_37
timestamp 1699142937
transform 1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_45
timestamp 1699142937
transform 1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_53
timestamp 1699142937
transform 1 0 5980 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_79
timestamp 1699142937
transform 1 0 8372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_3
timestamp 1699142937
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_11
timestamp 1699142937
transform 1 0 2116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_19
timestamp 1699142937
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_27
timestamp 1699142937
transform 1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_35
timestamp 1699142937
transform 1 0 4324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_43
timestamp 1699142937
transform 1 0 5060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1699142937
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1699142937
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_57
timestamp 1699142937
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1699142937
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_11
timestamp 1699142937
transform 1 0 2116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1699142937
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1699142937
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1699142937
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_37
timestamp 1699142937
transform 1 0 4508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_45
timestamp 1699142937
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_53
timestamp 1699142937
transform 1 0 5980 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_79
timestamp 1699142937
transform 1 0 8372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 1699142937
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_11
timestamp 1699142937
transform 1 0 2116 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_19
timestamp 1699142937
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_27
timestamp 1699142937
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_35
timestamp 1699142937
transform 1 0 4324 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_43
timestamp 1699142937
transform 1 0 5060 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1699142937
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1699142937
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_57
timestamp 1699142937
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_3
timestamp 1699142937
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_11
timestamp 1699142937
transform 1 0 2116 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_19
timestamp 1699142937
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1699142937
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_29
timestamp 1699142937
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_37
timestamp 1699142937
transform 1 0 4508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_45
timestamp 1699142937
transform 1 0 5244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_53
timestamp 1699142937
transform 1 0 5980 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_79
timestamp 1699142937
transform 1 0 8372 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1699142937
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_11
timestamp 1699142937
transform 1 0 2116 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_19
timestamp 1699142937
transform 1 0 2852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_27
timestamp 1699142937
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_35
timestamp 1699142937
transform 1 0 4324 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_43
timestamp 1699142937
transform 1 0 5060 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1699142937
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1699142937
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_57
timestamp 1699142937
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_3
timestamp 1699142937
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_11
timestamp 1699142937
transform 1 0 2116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_19
timestamp 1699142937
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1699142937
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_29
timestamp 1699142937
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_37
timestamp 1699142937
transform 1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_45
timestamp 1699142937
transform 1 0 5244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_53
timestamp 1699142937
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_61
timestamp 1699142937
transform 1 0 6716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_65
timestamp 1699142937
transform 1 0 7084 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 1699142937
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_11
timestamp 1699142937
transform 1 0 2116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_19
timestamp 1699142937
transform 1 0 2852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_27
timestamp 1699142937
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_35
timestamp 1699142937
transform 1 0 4324 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_43
timestamp 1699142937
transform 1 0 5060 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1699142937
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1699142937
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_57
timestamp 1699142937
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_79
timestamp 1699142937
transform 1 0 8372 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_3
timestamp 1699142937
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_11
timestamp 1699142937
transform 1 0 2116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_19
timestamp 1699142937
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1699142937
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_29
timestamp 1699142937
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_37
timestamp 1699142937
transform 1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_45
timestamp 1699142937
transform 1 0 5244 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_53
timestamp 1699142937
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_3
timestamp 1699142937
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_11
timestamp 1699142937
transform 1 0 2116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_19
timestamp 1699142937
transform 1 0 2852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_27
timestamp 1699142937
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_35
timestamp 1699142937
transform 1 0 4324 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_43
timestamp 1699142937
transform 1 0 5060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_49
timestamp 1699142937
transform 1 0 5612 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_80
timestamp 1699142937
transform 1 0 8464 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_3
timestamp 1699142937
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_11
timestamp 1699142937
transform 1 0 2116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_19
timestamp 1699142937
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1699142937
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_29
timestamp 1699142937
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_80
timestamp 1699142937
transform 1 0 8464 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_3
timestamp 1699142937
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_11
timestamp 1699142937
transform 1 0 2116 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_19
timestamp 1699142937
transform 1 0 2852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_27
timestamp 1699142937
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_35
timestamp 1699142937
transform 1 0 4324 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_43
timestamp 1699142937
transform 1 0 5060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1699142937
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1699142937
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_65
timestamp 1699142937
transform 1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_80
timestamp 1699142937
transform 1 0 8464 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_3
timestamp 1699142937
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_11
timestamp 1699142937
transform 1 0 2116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_19
timestamp 1699142937
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1699142937
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1699142937
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_37
timestamp 1699142937
transform 1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_45
timestamp 1699142937
transform 1 0 5244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_53
timestamp 1699142937
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_61
timestamp 1699142937
transform 1 0 6716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_69
timestamp 1699142937
transform 1 0 7452 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_3
timestamp 1699142937
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_11
timestamp 1699142937
transform 1 0 2116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_19
timestamp 1699142937
transform 1 0 2852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_27
timestamp 1699142937
transform 1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_35
timestamp 1699142937
transform 1 0 4324 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_57
timestamp 1699142937
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_61
timestamp 1699142937
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_74
timestamp 1699142937
transform 1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_3
timestamp 1699142937
transform 1 0 1380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_11
timestamp 1699142937
transform 1 0 2116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_19
timestamp 1699142937
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1699142937
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_29
timestamp 1699142937
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_37
timestamp 1699142937
transform 1 0 4508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_60
timestamp 1699142937
transform 1 0 6624 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_3
timestamp 1699142937
transform 1 0 1380 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_11
timestamp 1699142937
transform 1 0 2116 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_19
timestamp 1699142937
transform 1 0 2852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_27
timestamp 1699142937
transform 1 0 3588 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_35
timestamp 1699142937
transform 1 0 4324 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 1699142937
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_61
timestamp 1699142937
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_71
timestamp 1699142937
transform 1 0 7636 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_79
timestamp 1699142937
transform 1 0 8372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_3
timestamp 1699142937
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_11
timestamp 1699142937
transform 1 0 2116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_19
timestamp 1699142937
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1699142937
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_29
timestamp 1699142937
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_37
timestamp 1699142937
transform 1 0 4508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_45
timestamp 1699142937
transform 1 0 5244 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_57
timestamp 1699142937
transform 1 0 6348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_3
timestamp 1699142937
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_11
timestamp 1699142937
transform 1 0 2116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_19
timestamp 1699142937
transform 1 0 2852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_27
timestamp 1699142937
transform 1 0 3588 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_35
timestamp 1699142937
transform 1 0 4324 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_43
timestamp 1699142937
transform 1 0 5060 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_47
timestamp 1699142937
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1699142937
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_66
timestamp 1699142937
transform 1 0 7176 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_74
timestamp 1699142937
transform 1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_3
timestamp 1699142937
transform 1 0 1380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_11
timestamp 1699142937
transform 1 0 2116 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_19
timestamp 1699142937
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1699142937
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_29
timestamp 1699142937
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_37
timestamp 1699142937
transform 1 0 4508 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_60
timestamp 1699142937
transform 1 0 6624 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_76
timestamp 1699142937
transform 1 0 8096 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_3
timestamp 1699142937
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_11
timestamp 1699142937
transform 1 0 2116 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_19
timestamp 1699142937
transform 1 0 2852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_27
timestamp 1699142937
transform 1 0 3588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_35
timestamp 1699142937
transform 1 0 4324 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_43
timestamp 1699142937
transform 1 0 5060 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1699142937
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1699142937
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_57
timestamp 1699142937
transform 1 0 6348 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 1699142937
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_11
timestamp 1699142937
transform 1 0 2116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_19
timestamp 1699142937
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1699142937
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_29
timestamp 1699142937
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_37
timestamp 1699142937
transform 1 0 4508 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_57
timestamp 1699142937
transform 1 0 6348 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_70
timestamp 1699142937
transform 1 0 7544 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_78
timestamp 1699142937
transform 1 0 8280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_3
timestamp 1699142937
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_11
timestamp 1699142937
transform 1 0 2116 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_19
timestamp 1699142937
transform 1 0 2852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_27
timestamp 1699142937
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_35
timestamp 1699142937
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_57
timestamp 1699142937
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_3
timestamp 1699142937
transform 1 0 1380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_11
timestamp 1699142937
transform 1 0 2116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_19
timestamp 1699142937
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1699142937
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_29
timestamp 1699142937
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_37
timestamp 1699142937
transform 1 0 4508 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_45
timestamp 1699142937
transform 1 0 5244 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_53
timestamp 1699142937
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_61
timestamp 1699142937
transform 1 0 6716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_79
timestamp 1699142937
transform 1 0 8372 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_3
timestamp 1699142937
transform 1 0 1380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_11
timestamp 1699142937
transform 1 0 2116 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_19
timestamp 1699142937
transform 1 0 2852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_27
timestamp 1699142937
transform 1 0 3588 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_35
timestamp 1699142937
transform 1 0 4324 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_43
timestamp 1699142937
transform 1 0 5060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_57
timestamp 1699142937
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_79
timestamp 1699142937
transform 1 0 8372 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_3
timestamp 1699142937
transform 1 0 1380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_11
timestamp 1699142937
transform 1 0 2116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_19
timestamp 1699142937
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1699142937
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_29
timestamp 1699142937
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_37
timestamp 1699142937
transform 1 0 4508 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_60
timestamp 1699142937
transform 1 0 6624 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_3
timestamp 1699142937
transform 1 0 1380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_11
timestamp 1699142937
transform 1 0 2116 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_19
timestamp 1699142937
transform 1 0 2852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_27
timestamp 1699142937
transform 1 0 3588 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_35
timestamp 1699142937
transform 1 0 4324 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_52
timestamp 1699142937
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_57
timestamp 1699142937
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_61
timestamp 1699142937
transform 1 0 6716 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_73
timestamp 1699142937
transform 1 0 7820 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_3
timestamp 1699142937
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_11
timestamp 1699142937
transform 1 0 2116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_19
timestamp 1699142937
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1699142937
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_29
timestamp 1699142937
transform 1 0 3772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_37
timestamp 1699142937
transform 1 0 4508 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_3
timestamp 1699142937
transform 1 0 1380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_11
timestamp 1699142937
transform 1 0 2116 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_19
timestamp 1699142937
transform 1 0 2852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_27
timestamp 1699142937
transform 1 0 3588 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_35
timestamp 1699142937
transform 1 0 4324 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_46
timestamp 1699142937
transform 1 0 5336 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_57
timestamp 1699142937
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_65
timestamp 1699142937
transform 1 0 7084 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_73
timestamp 1699142937
transform 1 0 7820 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_3
timestamp 1699142937
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_11
timestamp 1699142937
transform 1 0 2116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_19
timestamp 1699142937
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1699142937
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_29
timestamp 1699142937
transform 1 0 3772 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_37
timestamp 1699142937
transform 1 0 4508 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_45
timestamp 1699142937
transform 1 0 5244 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_53
timestamp 1699142937
transform 1 0 5980 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_59
timestamp 1699142937
transform 1 0 6532 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_69
timestamp 1699142937
transform 1 0 7452 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_3
timestamp 1699142937
transform 1 0 1380 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_11
timestamp 1699142937
transform 1 0 2116 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_19
timestamp 1699142937
transform 1 0 2852 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_27
timestamp 1699142937
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_35
timestamp 1699142937
transform 1 0 4324 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_57
timestamp 1699142937
transform 1 0 6348 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_3
timestamp 1699142937
transform 1 0 1380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_11
timestamp 1699142937
transform 1 0 2116 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_19
timestamp 1699142937
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1699142937
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_29
timestamp 1699142937
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_37
timestamp 1699142937
transform 1 0 4508 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_55
timestamp 1699142937
transform 1 0 6164 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_70
timestamp 1699142937
transform 1 0 7544 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_78
timestamp 1699142937
transform 1 0 8280 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_3
timestamp 1699142937
transform 1 0 1380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_11
timestamp 1699142937
transform 1 0 2116 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_19
timestamp 1699142937
transform 1 0 2852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_27
timestamp 1699142937
transform 1 0 3588 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_35
timestamp 1699142937
transform 1 0 4324 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_46
timestamp 1699142937
transform 1 0 5336 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_57
timestamp 1699142937
transform 1 0 6348 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_3
timestamp 1699142937
transform 1 0 1380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_11
timestamp 1699142937
transform 1 0 2116 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_19
timestamp 1699142937
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1699142937
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_29
timestamp 1699142937
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_37
timestamp 1699142937
transform 1 0 4508 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_64
timestamp 1699142937
transform 1 0 6992 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_72
timestamp 1699142937
transform 1 0 7728 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_76
timestamp 1699142937
transform 1 0 8096 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_3
timestamp 1699142937
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_11
timestamp 1699142937
transform 1 0 2116 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_19
timestamp 1699142937
transform 1 0 2852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_27
timestamp 1699142937
transform 1 0 3588 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_35
timestamp 1699142937
transform 1 0 4324 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_43
timestamp 1699142937
transform 1 0 5060 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_57
timestamp 1699142937
transform 1 0 6348 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_73
timestamp 1699142937
transform 1 0 7820 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_3
timestamp 1699142937
transform 1 0 1380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_11
timestamp 1699142937
transform 1 0 2116 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_19
timestamp 1699142937
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1699142937
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_29
timestamp 1699142937
transform 1 0 3772 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_37
timestamp 1699142937
transform 1 0 4508 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_59
timestamp 1699142937
transform 1 0 6532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_3
timestamp 1699142937
transform 1 0 1380 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_11
timestamp 1699142937
transform 1 0 2116 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_19
timestamp 1699142937
transform 1 0 2852 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_27
timestamp 1699142937
transform 1 0 3588 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_35
timestamp 1699142937
transform 1 0 4324 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_43
timestamp 1699142937
transform 1 0 5060 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_54
timestamp 1699142937
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_70
timestamp 1699142937
transform 1 0 7544 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_78
timestamp 1699142937
transform 1 0 8280 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_3
timestamp 1699142937
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_11
timestamp 1699142937
transform 1 0 2116 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_19
timestamp 1699142937
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1699142937
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_29
timestamp 1699142937
transform 1 0 3772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_37
timestamp 1699142937
transform 1 0 4508 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_3
timestamp 1699142937
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_11
timestamp 1699142937
transform 1 0 2116 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_19
timestamp 1699142937
transform 1 0 2852 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_27
timestamp 1699142937
transform 1 0 3588 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_35
timestamp 1699142937
transform 1 0 4324 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_57
timestamp 1699142937
transform 1 0 6348 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_61
timestamp 1699142937
transform 1 0 6716 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_69
timestamp 1699142937
transform 1 0 7452 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_3
timestamp 1699142937
transform 1 0 1380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_11
timestamp 1699142937
transform 1 0 2116 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_19
timestamp 1699142937
transform 1 0 2852 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1699142937
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_29
timestamp 1699142937
transform 1 0 3772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_37
timestamp 1699142937
transform 1 0 4508 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_45
timestamp 1699142937
transform 1 0 5244 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_63
timestamp 1699142937
transform 1 0 6900 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_71
timestamp 1699142937
transform 1 0 7636 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_79
timestamp 1699142937
transform 1 0 8372 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_3
timestamp 1699142937
transform 1 0 1380 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_11
timestamp 1699142937
transform 1 0 2116 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_19
timestamp 1699142937
transform 1 0 2852 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_27
timestamp 1699142937
transform 1 0 3588 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_35
timestamp 1699142937
transform 1 0 4324 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_43
timestamp 1699142937
transform 1 0 5060 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_48
timestamp 1699142937
transform 1 0 5520 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_54
timestamp 1699142937
transform 1 0 6072 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_57
timestamp 1699142937
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_68
timestamp 1699142937
transform 1 0 7360 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_3
timestamp 1699142937
transform 1 0 1380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_11
timestamp 1699142937
transform 1 0 2116 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_19
timestamp 1699142937
transform 1 0 2852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1699142937
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_29
timestamp 1699142937
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_37
timestamp 1699142937
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_79
timestamp 1699142937
transform 1 0 8372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_3
timestamp 1699142937
transform 1 0 1380 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_11
timestamp 1699142937
transform 1 0 2116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_19
timestamp 1699142937
transform 1 0 2852 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_27
timestamp 1699142937
transform 1 0 3588 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_35
timestamp 1699142937
transform 1 0 4324 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_43
timestamp 1699142937
transform 1 0 5060 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1699142937
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_57
timestamp 1699142937
transform 1 0 6348 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_68
timestamp 1699142937
transform 1 0 7360 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_76
timestamp 1699142937
transform 1 0 8096 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_80
timestamp 1699142937
transform 1 0 8464 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_3
timestamp 1699142937
transform 1 0 1380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_11
timestamp 1699142937
transform 1 0 2116 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_19
timestamp 1699142937
transform 1 0 2852 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1699142937
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_29
timestamp 1699142937
transform 1 0 3772 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_37
timestamp 1699142937
transform 1 0 4508 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_61
timestamp 1699142937
transform 1 0 6716 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_69
timestamp 1699142937
transform 1 0 7452 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_77
timestamp 1699142937
transform 1 0 8188 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_3
timestamp 1699142937
transform 1 0 1380 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_11
timestamp 1699142937
transform 1 0 2116 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_19
timestamp 1699142937
transform 1 0 2852 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_27
timestamp 1699142937
transform 1 0 3588 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_35
timestamp 1699142937
transform 1 0 4324 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_43
timestamp 1699142937
transform 1 0 5060 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_47
timestamp 1699142937
transform 1 0 5428 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1699142937
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_57
timestamp 1699142937
transform 1 0 6348 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_63
timestamp 1699142937
transform 1 0 6900 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_67
timestamp 1699142937
transform 1 0 7268 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_75
timestamp 1699142937
transform 1 0 8004 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_3
timestamp 1699142937
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_11
timestamp 1699142937
transform 1 0 2116 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_19
timestamp 1699142937
transform 1 0 2852 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1699142937
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_29
timestamp 1699142937
transform 1 0 3772 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_37
timestamp 1699142937
transform 1 0 4508 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_48
timestamp 1699142937
transform 1 0 5520 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_56
timestamp 1699142937
transform 1 0 6256 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_60
timestamp 1699142937
transform 1 0 6624 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_3
timestamp 1699142937
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_11
timestamp 1699142937
transform 1 0 2116 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_19
timestamp 1699142937
transform 1 0 2852 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_27
timestamp 1699142937
transform 1 0 3588 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_57
timestamp 1699142937
transform 1 0 6348 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_78
timestamp 1699142937
transform 1 0 8280 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_3
timestamp 1699142937
transform 1 0 1380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_11
timestamp 1699142937
transform 1 0 2116 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_19
timestamp 1699142937
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1699142937
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_29
timestamp 1699142937
transform 1 0 3772 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_37
timestamp 1699142937
transform 1 0 4508 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_43
timestamp 1699142937
transform 1 0 5060 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_47
timestamp 1699142937
transform 1 0 5428 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_57
timestamp 1699142937
transform 1 0 6348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_3
timestamp 1699142937
transform 1 0 1380 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_11
timestamp 1699142937
transform 1 0 2116 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_19
timestamp 1699142937
transform 1 0 2852 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_27
timestamp 1699142937
transform 1 0 3588 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_35
timestamp 1699142937
transform 1 0 4324 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_57
timestamp 1699142937
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_61
timestamp 1699142937
transform 1 0 6716 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_71
timestamp 1699142937
transform 1 0 7636 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_3
timestamp 1699142937
transform 1 0 1380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_11
timestamp 1699142937
transform 1 0 2116 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_19
timestamp 1699142937
transform 1 0 2852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1699142937
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_29
timestamp 1699142937
transform 1 0 3772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_37
timestamp 1699142937
transform 1 0 4508 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82_45
timestamp 1699142937
transform 1 0 5244 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_71
timestamp 1699142937
transform 1 0 7636 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_3
timestamp 1699142937
transform 1 0 1380 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_11
timestamp 1699142937
transform 1 0 2116 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_19
timestamp 1699142937
transform 1 0 2852 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_27
timestamp 1699142937
transform 1 0 3588 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_35
timestamp 1699142937
transform 1 0 4324 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_57
timestamp 1699142937
transform 1 0 6348 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_3
timestamp 1699142937
transform 1 0 1380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_11
timestamp 1699142937
transform 1 0 2116 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_19
timestamp 1699142937
transform 1 0 2852 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 1699142937
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_29
timestamp 1699142937
transform 1 0 3772 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_37
timestamp 1699142937
transform 1 0 4508 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_43
timestamp 1699142937
transform 1 0 5060 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_56
timestamp 1699142937
transform 1 0 6256 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_71
timestamp 1699142937
transform 1 0 7636 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_84_79
timestamp 1699142937
transform 1 0 8372 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_3
timestamp 1699142937
transform 1 0 1380 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_11
timestamp 1699142937
transform 1 0 2116 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_19
timestamp 1699142937
transform 1 0 2852 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_27
timestamp 1699142937
transform 1 0 3588 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_35
timestamp 1699142937
transform 1 0 4324 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_46
timestamp 1699142937
transform 1 0 5336 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_57
timestamp 1699142937
transform 1 0 6348 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_3
timestamp 1699142937
transform 1 0 1380 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_11
timestamp 1699142937
transform 1 0 2116 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_19
timestamp 1699142937
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1699142937
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_29
timestamp 1699142937
transform 1 0 3772 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_86_37
timestamp 1699142937
transform 1 0 4508 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_59
timestamp 1699142937
transform 1 0 6532 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_86_72
timestamp 1699142937
transform 1 0 7728 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_76
timestamp 1699142937
transform 1 0 8096 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_3
timestamp 1699142937
transform 1 0 1380 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_11
timestamp 1699142937
transform 1 0 2116 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_19
timestamp 1699142937
transform 1 0 2852 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_27
timestamp 1699142937
transform 1 0 3588 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87_35
timestamp 1699142937
transform 1 0 4324 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_48
timestamp 1699142937
transform 1 0 5520 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87_57
timestamp 1699142937
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_70
timestamp 1699142937
transform 1 0 7544 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_76
timestamp 1699142937
transform 1 0 8096 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_3
timestamp 1699142937
transform 1 0 1380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_11
timestamp 1699142937
transform 1 0 2116 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_19
timestamp 1699142937
transform 1 0 2852 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 1699142937
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_29
timestamp 1699142937
transform 1 0 3772 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_57
timestamp 1699142937
transform 1 0 6348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_3
timestamp 1699142937
transform 1 0 1380 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_11
timestamp 1699142937
transform 1 0 2116 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_19
timestamp 1699142937
transform 1 0 2852 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_27
timestamp 1699142937
transform 1 0 3588 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_35
timestamp 1699142937
transform 1 0 4324 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_41
timestamp 1699142937
transform 1 0 4876 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_45
timestamp 1699142937
transform 1 0 5244 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 1699142937
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_89_57
timestamp 1699142937
transform 1 0 6348 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_69
timestamp 1699142937
transform 1 0 7452 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_77
timestamp 1699142937
transform 1 0 8188 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_3
timestamp 1699142937
transform 1 0 1380 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_11
timestamp 1699142937
transform 1 0 2116 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_19
timestamp 1699142937
transform 1 0 2852 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 1699142937
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_29
timestamp 1699142937
transform 1 0 3772 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90_37
timestamp 1699142937
transform 1 0 4508 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_44
timestamp 1699142937
transform 1 0 5152 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90_54
timestamp 1699142937
transform 1 0 6072 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_3
timestamp 1699142937
transform 1 0 1380 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_11
timestamp 1699142937
transform 1 0 2116 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_19
timestamp 1699142937
transform 1 0 2852 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_27
timestamp 1699142937
transform 1 0 3588 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_35
timestamp 1699142937
transform 1 0 4324 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_57
timestamp 1699142937
transform 1 0 6348 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_65
timestamp 1699142937
transform 1 0 7084 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_73
timestamp 1699142937
transform 1 0 7820 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_3
timestamp 1699142937
transform 1 0 1380 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_11
timestamp 1699142937
transform 1 0 2116 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_19
timestamp 1699142937
transform 1 0 2852 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1699142937
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_29
timestamp 1699142937
transform 1 0 3772 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_37
timestamp 1699142937
transform 1 0 4508 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_45
timestamp 1699142937
transform 1 0 5244 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_53
timestamp 1699142937
transform 1 0 5980 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_59
timestamp 1699142937
transform 1 0 6532 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_69
timestamp 1699142937
transform 1 0 7452 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_3
timestamp 1699142937
transform 1 0 1380 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_11
timestamp 1699142937
transform 1 0 2116 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_19
timestamp 1699142937
transform 1 0 2852 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_27
timestamp 1699142937
transform 1 0 3588 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_35
timestamp 1699142937
transform 1 0 4324 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_57
timestamp 1699142937
transform 1 0 6348 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_3
timestamp 1699142937
transform 1 0 1380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_11
timestamp 1699142937
transform 1 0 2116 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_19
timestamp 1699142937
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1699142937
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_29
timestamp 1699142937
transform 1 0 3772 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_37
timestamp 1699142937
transform 1 0 4508 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_41
timestamp 1699142937
transform 1 0 4876 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_54
timestamp 1699142937
transform 1 0 6072 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_69
timestamp 1699142937
transform 1 0 7452 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_77
timestamp 1699142937
transform 1 0 8188 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_3
timestamp 1699142937
transform 1 0 1380 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_11
timestamp 1699142937
transform 1 0 2116 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_19
timestamp 1699142937
transform 1 0 2852 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_27
timestamp 1699142937
transform 1 0 3588 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_35
timestamp 1699142937
transform 1 0 4324 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_41
timestamp 1699142937
transform 1 0 4876 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_54
timestamp 1699142937
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_57
timestamp 1699142937
transform 1 0 6348 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_3
timestamp 1699142937
transform 1 0 1380 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_11
timestamp 1699142937
transform 1 0 2116 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_19
timestamp 1699142937
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1699142937
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_29
timestamp 1699142937
transform 1 0 3772 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_57
timestamp 1699142937
transform 1 0 6348 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96_65
timestamp 1699142937
transform 1 0 7084 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_73
timestamp 1699142937
transform 1 0 7820 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_3
timestamp 1699142937
transform 1 0 1380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_11
timestamp 1699142937
transform 1 0 2116 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_19
timestamp 1699142937
transform 1 0 2852 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_27
timestamp 1699142937
transform 1 0 3588 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_35
timestamp 1699142937
transform 1 0 4324 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_43
timestamp 1699142937
transform 1 0 5060 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 1699142937
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 1699142937
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_57
timestamp 1699142937
transform 1 0 6348 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_69
timestamp 1699142937
transform 1 0 7452 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_3
timestamp 1699142937
transform 1 0 1380 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_11
timestamp 1699142937
transform 1 0 2116 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_19
timestamp 1699142937
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1699142937
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_29
timestamp 1699142937
transform 1 0 3772 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_57
timestamp 1699142937
transform 1 0 6348 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_3
timestamp 1699142937
transform 1 0 1380 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_11
timestamp 1699142937
transform 1 0 2116 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_19
timestamp 1699142937
transform 1 0 2852 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_27
timestamp 1699142937
transform 1 0 3588 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_35
timestamp 1699142937
transform 1 0 4324 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_41
timestamp 1699142937
transform 1 0 4876 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_54
timestamp 1699142937
transform 1 0 6072 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_70
timestamp 1699142937
transform 1 0 7544 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_99_78
timestamp 1699142937
transform 1 0 8280 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_3
timestamp 1699142937
transform 1 0 1380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_11
timestamp 1699142937
transform 1 0 2116 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_19
timestamp 1699142937
transform 1 0 2852 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 1699142937
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_29
timestamp 1699142937
transform 1 0 3772 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_37
timestamp 1699142937
transform 1 0 4508 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_60
timestamp 1699142937
transform 1 0 6624 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_3
timestamp 1699142937
transform 1 0 1380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_11
timestamp 1699142937
transform 1 0 2116 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_19
timestamp 1699142937
transform 1 0 2852 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_27
timestamp 1699142937
transform 1 0 3588 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_35
timestamp 1699142937
transform 1 0 4324 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_57
timestamp 1699142937
transform 1 0 6348 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_61
timestamp 1699142937
transform 1 0 6716 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_65
timestamp 1699142937
transform 1 0 7084 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_77
timestamp 1699142937
transform 1 0 8188 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_3
timestamp 1699142937
transform 1 0 1380 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_11
timestamp 1699142937
transform 1 0 2116 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_19
timestamp 1699142937
transform 1 0 2852 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_27
timestamp 1699142937
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_29
timestamp 1699142937
transform 1 0 3772 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_37
timestamp 1699142937
transform 1 0 4508 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_41
timestamp 1699142937
transform 1 0 4876 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_45
timestamp 1699142937
transform 1 0 5244 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_53
timestamp 1699142937
transform 1 0 5980 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_70
timestamp 1699142937
transform 1 0 7544 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_74
timestamp 1699142937
transform 1 0 7912 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_3
timestamp 1699142937
transform 1 0 1380 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_11
timestamp 1699142937
transform 1 0 2116 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_19
timestamp 1699142937
transform 1 0 2852 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_27
timestamp 1699142937
transform 1 0 3588 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_35
timestamp 1699142937
transform 1 0 4324 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_57
timestamp 1699142937
transform 1 0 6348 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_3
timestamp 1699142937
transform 1 0 1380 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_11
timestamp 1699142937
transform 1 0 2116 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_19
timestamp 1699142937
transform 1 0 2852 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_27
timestamp 1699142937
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_29
timestamp 1699142937
transform 1 0 3772 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_37
timestamp 1699142937
transform 1 0 4508 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_54
timestamp 1699142937
transform 1 0 6072 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_60
timestamp 1699142937
transform 1 0 6624 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_70
timestamp 1699142937
transform 1 0 7544 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_74
timestamp 1699142937
transform 1 0 7912 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_3
timestamp 1699142937
transform 1 0 1380 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_11
timestamp 1699142937
transform 1 0 2116 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_19
timestamp 1699142937
transform 1 0 2852 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_27
timestamp 1699142937
transform 1 0 3588 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_35
timestamp 1699142937
transform 1 0 4324 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_57
timestamp 1699142937
transform 1 0 6348 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_3
timestamp 1699142937
transform 1 0 1380 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_11
timestamp 1699142937
transform 1 0 2116 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_19
timestamp 1699142937
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_27
timestamp 1699142937
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_29
timestamp 1699142937
transform 1 0 3772 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106_37
timestamp 1699142937
transform 1 0 4508 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_53
timestamp 1699142937
transform 1 0 5980 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_59
timestamp 1699142937
transform 1 0 6532 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_69
timestamp 1699142937
transform 1 0 7452 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_3
timestamp 1699142937
transform 1 0 1380 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_11
timestamp 1699142937
transform 1 0 2116 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_19
timestamp 1699142937
transform 1 0 2852 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_27
timestamp 1699142937
transform 1 0 3588 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_35
timestamp 1699142937
transform 1 0 4324 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_39
timestamp 1699142937
transform 1 0 4692 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_43
timestamp 1699142937
transform 1 0 5060 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107_53
timestamp 1699142937
transform 1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_57
timestamp 1699142937
transform 1 0 6348 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_3
timestamp 1699142937
transform 1 0 1380 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_11
timestamp 1699142937
transform 1 0 2116 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_19
timestamp 1699142937
transform 1 0 2852 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_27
timestamp 1699142937
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_29
timestamp 1699142937
transform 1 0 3772 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_35
timestamp 1699142937
transform 1 0 4324 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_56
timestamp 1699142937
transform 1 0 6256 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_71
timestamp 1699142937
transform 1 0 7636 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_3
timestamp 1699142937
transform 1 0 1380 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_11
timestamp 1699142937
transform 1 0 2116 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_19
timestamp 1699142937
transform 1 0 2852 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_27
timestamp 1699142937
transform 1 0 3588 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_35
timestamp 1699142937
transform 1 0 4324 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_43
timestamp 1699142937
transform 1 0 5060 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_51
timestamp 1699142937
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_55
timestamp 1699142937
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_57
timestamp 1699142937
transform 1 0 6348 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_70
timestamp 1699142937
transform 1 0 7544 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109_78
timestamp 1699142937
transform 1 0 8280 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_3
timestamp 1699142937
transform 1 0 1380 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_11
timestamp 1699142937
transform 1 0 2116 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_19
timestamp 1699142937
transform 1 0 2852 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_27
timestamp 1699142937
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_29
timestamp 1699142937
transform 1 0 3772 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_110_55
timestamp 1699142937
transform 1 0 6164 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_3
timestamp 1699142937
transform 1 0 1380 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_11
timestamp 1699142937
transform 1 0 2116 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_19
timestamp 1699142937
transform 1 0 2852 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_27
timestamp 1699142937
transform 1 0 3588 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_35
timestamp 1699142937
transform 1 0 4324 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_39
timestamp 1699142937
transform 1 0 4692 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_43
timestamp 1699142937
transform 1 0 5060 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_111_53
timestamp 1699142937
transform 1 0 5980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_57
timestamp 1699142937
transform 1 0 6348 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_65
timestamp 1699142937
transform 1 0 7084 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_73
timestamp 1699142937
transform 1 0 7820 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_3
timestamp 1699142937
transform 1 0 1380 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_11
timestamp 1699142937
transform 1 0 2116 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_19
timestamp 1699142937
transform 1 0 2852 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_27
timestamp 1699142937
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_29
timestamp 1699142937
transform 1 0 3772 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112_55
timestamp 1699142937
transform 1 0 6164 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_3
timestamp 1699142937
transform 1 0 1380 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_11
timestamp 1699142937
transform 1 0 2116 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_19
timestamp 1699142937
transform 1 0 2852 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113_27
timestamp 1699142937
transform 1 0 3588 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_35
timestamp 1699142937
transform 1 0 4324 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_39
timestamp 1699142937
transform 1 0 4692 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113_43
timestamp 1699142937
transform 1 0 5060 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113_54
timestamp 1699142937
transform 1 0 6072 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_57
timestamp 1699142937
transform 1 0 6348 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113_78
timestamp 1699142937
transform 1 0 8280 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_3
timestamp 1699142937
transform 1 0 1380 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_11
timestamp 1699142937
transform 1 0 2116 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_19
timestamp 1699142937
transform 1 0 2852 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_27
timestamp 1699142937
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_29
timestamp 1699142937
transform 1 0 3772 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_37
timestamp 1699142937
transform 1 0 4508 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_45
timestamp 1699142937
transform 1 0 5244 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_53
timestamp 1699142937
transform 1 0 5980 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_57
timestamp 1699142937
transform 1 0 6348 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_3
timestamp 1699142937
transform 1 0 1380 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_11
timestamp 1699142937
transform 1 0 2116 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_19
timestamp 1699142937
transform 1 0 2852 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_27
timestamp 1699142937
transform 1 0 3588 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_115_35
timestamp 1699142937
transform 1 0 4324 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_52
timestamp 1699142937
transform 1 0 5888 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_57
timestamp 1699142937
transform 1 0 6348 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_61
timestamp 1699142937
transform 1 0 6716 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_115_65
timestamp 1699142937
transform 1 0 7084 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_73
timestamp 1699142937
transform 1 0 7820 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_3
timestamp 1699142937
transform 1 0 1380 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_11
timestamp 1699142937
transform 1 0 2116 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_19
timestamp 1699142937
transform 1 0 2852 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_27
timestamp 1699142937
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_29
timestamp 1699142937
transform 1 0 3772 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116_37
timestamp 1699142937
transform 1 0 4508 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_72
timestamp 1699142937
transform 1 0 7728 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_76
timestamp 1699142937
transform 1 0 8096 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_3
timestamp 1699142937
transform 1 0 1380 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_11
timestamp 1699142937
transform 1 0 2116 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_19
timestamp 1699142937
transform 1 0 2852 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_27
timestamp 1699142937
transform 1 0 3588 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_35
timestamp 1699142937
transform 1 0 4324 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117_43
timestamp 1699142937
transform 1 0 5060 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117_48
timestamp 1699142937
transform 1 0 5520 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_57
timestamp 1699142937
transform 1 0 6348 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_3
timestamp 1699142937
transform 1 0 1380 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_11
timestamp 1699142937
transform 1 0 2116 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_19
timestamp 1699142937
transform 1 0 2852 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_27
timestamp 1699142937
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_29
timestamp 1699142937
transform 1 0 3772 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_118_37
timestamp 1699142937
transform 1 0 4508 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_80
timestamp 1699142937
transform 1 0 8464 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_3
timestamp 1699142937
transform 1 0 1380 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_11
timestamp 1699142937
transform 1 0 2116 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_19
timestamp 1699142937
transform 1 0 2852 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_27
timestamp 1699142937
transform 1 0 3588 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_35
timestamp 1699142937
transform 1 0 4324 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_43
timestamp 1699142937
transform 1 0 5060 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_51
timestamp 1699142937
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_55
timestamp 1699142937
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_69
timestamp 1699142937
transform 1 0 7452 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_3
timestamp 1699142937
transform 1 0 1380 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_11
timestamp 1699142937
transform 1 0 2116 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_19
timestamp 1699142937
transform 1 0 2852 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_27
timestamp 1699142937
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_29
timestamp 1699142937
transform 1 0 3772 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_120_37
timestamp 1699142937
transform 1 0 4508 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_60
timestamp 1699142937
transform 1 0 6624 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_3
timestamp 1699142937
transform 1 0 1380 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_11
timestamp 1699142937
transform 1 0 2116 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_19
timestamp 1699142937
transform 1 0 2852 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_27
timestamp 1699142937
transform 1 0 3588 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_35
timestamp 1699142937
transform 1 0 4324 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_43
timestamp 1699142937
transform 1 0 5060 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_57
timestamp 1699142937
transform 1 0 6348 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_61
timestamp 1699142937
transform 1 0 6716 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_71
timestamp 1699142937
transform 1 0 7636 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_3
timestamp 1699142937
transform 1 0 1380 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_11
timestamp 1699142937
transform 1 0 2116 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_19
timestamp 1699142937
transform 1 0 2852 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_27
timestamp 1699142937
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_29
timestamp 1699142937
transform 1 0 3772 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_37
timestamp 1699142937
transform 1 0 4508 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_43
timestamp 1699142937
transform 1 0 5060 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_47
timestamp 1699142937
transform 1 0 5428 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_57
timestamp 1699142937
transform 1 0 6348 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_3
timestamp 1699142937
transform 1 0 1380 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_11
timestamp 1699142937
transform 1 0 2116 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_19
timestamp 1699142937
transform 1 0 2852 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_27
timestamp 1699142937
transform 1 0 3588 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_35
timestamp 1699142937
transform 1 0 4324 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123_57
timestamp 1699142937
transform 1 0 6348 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_61
timestamp 1699142937
transform 1 0 6716 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_71
timestamp 1699142937
transform 1 0 7636 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_3
timestamp 1699142937
transform 1 0 1380 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_11
timestamp 1699142937
transform 1 0 2116 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_19
timestamp 1699142937
transform 1 0 2852 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_27
timestamp 1699142937
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_29
timestamp 1699142937
transform 1 0 3772 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_37
timestamp 1699142937
transform 1 0 4508 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_45
timestamp 1699142937
transform 1 0 5244 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_53
timestamp 1699142937
transform 1 0 5980 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124_61
timestamp 1699142937
transform 1 0 6716 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_124_72
timestamp 1699142937
transform 1 0 7728 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_80
timestamp 1699142937
transform 1 0 8464 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_3
timestamp 1699142937
transform 1 0 1380 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_11
timestamp 1699142937
transform 1 0 2116 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_19
timestamp 1699142937
transform 1 0 2852 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125_27
timestamp 1699142937
transform 1 0 3588 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_35
timestamp 1699142937
transform 1 0 4324 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125_57
timestamp 1699142937
transform 1 0 6348 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126_3
timestamp 1699142937
transform 1 0 1380 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126_11
timestamp 1699142937
transform 1 0 2116 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126_19
timestamp 1699142937
transform 1 0 2852 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_27
timestamp 1699142937
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126_29
timestamp 1699142937
transform 1 0 3772 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_126_37
timestamp 1699142937
transform 1 0 4508 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_43
timestamp 1699142937
transform 1 0 5060 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_47
timestamp 1699142937
transform 1 0 5428 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_126_57
timestamp 1699142937
transform 1 0 6348 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_63
timestamp 1699142937
transform 1 0 6900 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126_67
timestamp 1699142937
transform 1 0 7268 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126_75
timestamp 1699142937
transform 1 0 8004 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_3
timestamp 1699142937
transform 1 0 1380 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_11
timestamp 1699142937
transform 1 0 2116 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_19
timestamp 1699142937
transform 1 0 2852 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_27
timestamp 1699142937
transform 1 0 3588 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_35
timestamp 1699142937
transform 1 0 4324 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127_43
timestamp 1699142937
transform 1 0 5060 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127_48
timestamp 1699142937
transform 1 0 5520 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_128_3
timestamp 1699142937
transform 1 0 1380 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_128_11
timestamp 1699142937
transform 1 0 2116 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_128_19
timestamp 1699142937
transform 1 0 2852 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_27
timestamp 1699142937
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_128_29
timestamp 1699142937
transform 1 0 3772 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128_37
timestamp 1699142937
transform 1 0 4508 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_60
timestamp 1699142937
transform 1 0 6624 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_3
timestamp 1699142937
transform 1 0 1380 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_11
timestamp 1699142937
transform 1 0 2116 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_19
timestamp 1699142937
transform 1 0 2852 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_27
timestamp 1699142937
transform 1 0 3588 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_35
timestamp 1699142937
transform 1 0 4324 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129_43
timestamp 1699142937
transform 1 0 5060 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_129_50
timestamp 1699142937
transform 1 0 5704 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129_69
timestamp 1699142937
transform 1 0 7452 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129_77
timestamp 1699142937
transform 1 0 8188 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130_3
timestamp 1699142937
transform 1 0 1380 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130_11
timestamp 1699142937
transform 1 0 2116 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130_19
timestamp 1699142937
transform 1 0 2852 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_27
timestamp 1699142937
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130_29
timestamp 1699142937
transform 1 0 3772 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_130_37
timestamp 1699142937
transform 1 0 4508 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_3
timestamp 1699142937
transform 1 0 1380 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_11
timestamp 1699142937
transform 1 0 2116 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_19
timestamp 1699142937
transform 1 0 2852 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_27
timestamp 1699142937
transform 1 0 3588 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_35
timestamp 1699142937
transform 1 0 4324 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131_43
timestamp 1699142937
transform 1 0 5060 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131_51
timestamp 1699142937
transform 1 0 5796 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_55
timestamp 1699142937
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_3
timestamp 1699142937
transform 1 0 1380 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_11
timestamp 1699142937
transform 1 0 2116 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_19
timestamp 1699142937
transform 1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_27
timestamp 1699142937
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_29
timestamp 1699142937
transform 1 0 3772 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_37
timestamp 1699142937
transform 1 0 4508 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_45
timestamp 1699142937
transform 1 0 5244 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_53
timestamp 1699142937
transform 1 0 5980 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_61
timestamp 1699142937
transform 1 0 6716 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_69
timestamp 1699142937
transform 1 0 7452 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_3
timestamp 1699142937
transform 1 0 1380 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_11
timestamp 1699142937
transform 1 0 2116 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_19
timestamp 1699142937
transform 1 0 2852 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_27
timestamp 1699142937
transform 1 0 3588 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_35
timestamp 1699142937
transform 1 0 4324 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_43
timestamp 1699142937
transform 1 0 5060 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133_51
timestamp 1699142937
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_55
timestamp 1699142937
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_57
timestamp 1699142937
transform 1 0 6348 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_65
timestamp 1699142937
transform 1 0 7084 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133_73
timestamp 1699142937
transform 1 0 7820 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_3
timestamp 1699142937
transform 1 0 1380 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_11
timestamp 1699142937
transform 1 0 2116 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_19
timestamp 1699142937
transform 1 0 2852 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_27
timestamp 1699142937
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_29
timestamp 1699142937
transform 1 0 3772 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_37
timestamp 1699142937
transform 1 0 4508 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_45
timestamp 1699142937
transform 1 0 5244 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_53
timestamp 1699142937
transform 1 0 5980 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_61
timestamp 1699142937
transform 1 0 6716 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_69
timestamp 1699142937
transform 1 0 7452 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134_77
timestamp 1699142937
transform 1 0 8188 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_3
timestamp 1699142937
transform 1 0 1380 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_11
timestamp 1699142937
transform 1 0 2116 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_19
timestamp 1699142937
transform 1 0 2852 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_27
timestamp 1699142937
transform 1 0 3588 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_35
timestamp 1699142937
transform 1 0 4324 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_43
timestamp 1699142937
transform 1 0 5060 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135_51
timestamp 1699142937
transform 1 0 5796 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_55
timestamp 1699142937
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_57
timestamp 1699142937
transform 1 0 6348 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_65
timestamp 1699142937
transform 1 0 7084 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135_73
timestamp 1699142937
transform 1 0 7820 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_3
timestamp 1699142937
transform 1 0 1380 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_11
timestamp 1699142937
transform 1 0 2116 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_19
timestamp 1699142937
transform 1 0 2852 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_27
timestamp 1699142937
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_29
timestamp 1699142937
transform 1 0 3772 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_37
timestamp 1699142937
transform 1 0 4508 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_45
timestamp 1699142937
transform 1 0 5244 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_53
timestamp 1699142937
transform 1 0 5980 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_61
timestamp 1699142937
transform 1 0 6716 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_69
timestamp 1699142937
transform 1 0 7452 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136_77
timestamp 1699142937
transform 1 0 8188 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_3
timestamp 1699142937
transform 1 0 1380 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_11
timestamp 1699142937
transform 1 0 2116 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_19
timestamp 1699142937
transform 1 0 2852 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_27
timestamp 1699142937
transform 1 0 3588 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_35
timestamp 1699142937
transform 1 0 4324 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_43
timestamp 1699142937
transform 1 0 5060 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_137_51
timestamp 1699142937
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_55
timestamp 1699142937
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_57
timestamp 1699142937
transform 1 0 6348 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_65
timestamp 1699142937
transform 1 0 7084 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137_73
timestamp 1699142937
transform 1 0 7820 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_3
timestamp 1699142937
transform 1 0 1380 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_138_11
timestamp 1699142937
transform 1 0 2116 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_15
timestamp 1699142937
transform 1 0 2484 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_20
timestamp 1699142937
transform 1 0 2944 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_29
timestamp 1699142937
transform 1 0 3772 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_37
timestamp 1699142937
transform 1 0 4508 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_45
timestamp 1699142937
transform 1 0 5244 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_138_53
timestamp 1699142937
transform 1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_57
timestamp 1699142937
transform 1 0 6348 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_65
timestamp 1699142937
transform 1 0 7084 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_73
timestamp 1699142937
transform 1 0 7820 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1699142937
transform -1 0 6164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1699142937
transform -1 0 7084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1699142937
transform 1 0 7084 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1699142937
transform 1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1699142937
transform 1 0 7084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1699142937
transform 1 0 6992 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1699142937
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1699142937
transform 1 0 7084 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1699142937
transform -1 0 8556 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1699142937
transform -1 0 8556 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1699142937
transform -1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1699142937
transform -1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1699142937
transform 1 0 6532 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1699142937
transform 1 0 6992 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1699142937
transform 1 0 6992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1699142937
transform -1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1699142937
transform -1 0 8464 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1699142937
transform -1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1699142937
transform -1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1699142937
transform -1 0 8556 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1699142937
transform -1 0 7728 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1699142937
transform 1 0 8280 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1699142937
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1699142937
transform -1 0 6808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1699142937
transform -1 0 6992 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1699142937
transform -1 0 7176 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1699142937
transform -1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1699142937
transform 1 0 8004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1699142937
transform 1 0 8280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1699142937
transform -1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1699142937
transform -1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1699142937
transform -1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1699142937
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1699142937
transform -1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1699142937
transform 1 0 8280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1699142937
transform -1 0 6808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1699142937
transform -1 0 7360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1699142937
transform -1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1699142937
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1699142937
transform -1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1699142937
transform 1 0 2576 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1699142937
transform -1 0 7820 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1699142937
transform 1 0 8188 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1699142937
transform 1 0 8188 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1699142937
transform 1 0 8188 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1699142937
transform 1 0 8188 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1699142937
transform 1 0 8004 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1699142937
transform 1 0 8188 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1699142937
transform 1 0 8188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1699142937
transform 1 0 8188 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1699142937
transform 1 0 8188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1699142937
transform 1 0 8188 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1699142937
transform 1 0 8188 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1699142937
transform 1 0 8188 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1699142937
transform 1 0 8188 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1699142937
transform 1 0 8188 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1699142937
transform 1 0 7820 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1699142937
transform 1 0 8188 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1699142937
transform 1 0 8004 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1699142937
transform 1 0 8188 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1699142937
transform 1 0 8188 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1699142937
transform 1 0 8188 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1699142937
transform 1 0 8004 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1699142937
transform 1 0 8188 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1699142937
transform 1 0 8188 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1699142937
transform 1 0 8188 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1699142937
transform 1 0 8188 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1699142937
transform 1 0 8188 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1699142937
transform 1 0 8188 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1699142937
transform 1 0 8188 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1699142937
transform 1 0 8188 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output52
timestamp 1699142937
transform -1 0 7820 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output53
timestamp 1699142937
transform 1 0 7636 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 1699142937
transform 1 0 8004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1699142937
transform -1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_139
timestamp 1699142937
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1699142937
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_140
timestamp 1699142937
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1699142937
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_141
timestamp 1699142937
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1699142937
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_142
timestamp 1699142937
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1699142937
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_143
timestamp 1699142937
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1699142937
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_144
timestamp 1699142937
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1699142937
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_145
timestamp 1699142937
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1699142937
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_146
timestamp 1699142937
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1699142937
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_147
timestamp 1699142937
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1699142937
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_148
timestamp 1699142937
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1699142937
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_149
timestamp 1699142937
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1699142937
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_150
timestamp 1699142937
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1699142937
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_151
timestamp 1699142937
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1699142937
transform -1 0 8832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_152
timestamp 1699142937
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1699142937
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_153
timestamp 1699142937
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1699142937
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_154
timestamp 1699142937
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1699142937
transform -1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_155
timestamp 1699142937
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1699142937
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_156
timestamp 1699142937
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1699142937
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_157
timestamp 1699142937
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1699142937
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_158
timestamp 1699142937
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1699142937
transform -1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_159
timestamp 1699142937
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1699142937
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_160
timestamp 1699142937
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1699142937
transform -1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_161
timestamp 1699142937
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1699142937
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_162
timestamp 1699142937
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1699142937
transform -1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_163
timestamp 1699142937
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1699142937
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_164
timestamp 1699142937
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1699142937
transform -1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_165
timestamp 1699142937
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1699142937
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_166
timestamp 1699142937
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1699142937
transform -1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_167
timestamp 1699142937
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1699142937
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_168
timestamp 1699142937
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1699142937
transform -1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_169
timestamp 1699142937
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1699142937
transform -1 0 8832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_170
timestamp 1699142937
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1699142937
transform -1 0 8832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_171
timestamp 1699142937
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1699142937
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_172
timestamp 1699142937
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1699142937
transform -1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_173
timestamp 1699142937
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1699142937
transform -1 0 8832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_174
timestamp 1699142937
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1699142937
transform -1 0 8832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_175
timestamp 1699142937
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1699142937
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_176
timestamp 1699142937
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1699142937
transform -1 0 8832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_177
timestamp 1699142937
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1699142937
transform -1 0 8832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_178
timestamp 1699142937
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1699142937
transform -1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_179
timestamp 1699142937
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1699142937
transform -1 0 8832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_180
timestamp 1699142937
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1699142937
transform -1 0 8832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_181
timestamp 1699142937
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1699142937
transform -1 0 8832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_182
timestamp 1699142937
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1699142937
transform -1 0 8832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_183
timestamp 1699142937
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1699142937
transform -1 0 8832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_184
timestamp 1699142937
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1699142937
transform -1 0 8832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_185
timestamp 1699142937
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1699142937
transform -1 0 8832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_186
timestamp 1699142937
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1699142937
transform -1 0 8832 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_187
timestamp 1699142937
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1699142937
transform -1 0 8832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_188
timestamp 1699142937
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1699142937
transform -1 0 8832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_189
timestamp 1699142937
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1699142937
transform -1 0 8832 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_190
timestamp 1699142937
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1699142937
transform -1 0 8832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_191
timestamp 1699142937
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1699142937
transform -1 0 8832 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_192
timestamp 1699142937
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1699142937
transform -1 0 8832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_193
timestamp 1699142937
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1699142937
transform -1 0 8832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_194
timestamp 1699142937
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1699142937
transform -1 0 8832 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_195
timestamp 1699142937
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1699142937
transform -1 0 8832 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_196
timestamp 1699142937
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1699142937
transform -1 0 8832 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_197
timestamp 1699142937
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1699142937
transform -1 0 8832 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_198
timestamp 1699142937
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1699142937
transform -1 0 8832 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_199
timestamp 1699142937
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1699142937
transform -1 0 8832 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_200
timestamp 1699142937
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1699142937
transform -1 0 8832 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_201
timestamp 1699142937
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1699142937
transform -1 0 8832 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_202
timestamp 1699142937
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1699142937
transform -1 0 8832 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_203
timestamp 1699142937
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1699142937
transform -1 0 8832 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_204
timestamp 1699142937
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1699142937
transform -1 0 8832 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_205
timestamp 1699142937
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1699142937
transform -1 0 8832 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_206
timestamp 1699142937
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1699142937
transform -1 0 8832 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_207
timestamp 1699142937
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1699142937
transform -1 0 8832 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_208
timestamp 1699142937
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1699142937
transform -1 0 8832 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_209
timestamp 1699142937
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1699142937
transform -1 0 8832 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_210
timestamp 1699142937
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1699142937
transform -1 0 8832 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_211
timestamp 1699142937
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1699142937
transform -1 0 8832 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_212
timestamp 1699142937
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1699142937
transform -1 0 8832 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_213
timestamp 1699142937
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1699142937
transform -1 0 8832 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_214
timestamp 1699142937
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1699142937
transform -1 0 8832 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_215
timestamp 1699142937
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1699142937
transform -1 0 8832 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_216
timestamp 1699142937
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1699142937
transform -1 0 8832 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_217
timestamp 1699142937
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1699142937
transform -1 0 8832 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_218
timestamp 1699142937
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1699142937
transform -1 0 8832 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_219
timestamp 1699142937
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1699142937
transform -1 0 8832 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_220
timestamp 1699142937
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 1699142937
transform -1 0 8832 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_221
timestamp 1699142937
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 1699142937
transform -1 0 8832 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_222
timestamp 1699142937
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 1699142937
transform -1 0 8832 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_223
timestamp 1699142937
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 1699142937
transform -1 0 8832 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_224
timestamp 1699142937
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 1699142937
transform -1 0 8832 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_225
timestamp 1699142937
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 1699142937
transform -1 0 8832 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_226
timestamp 1699142937
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 1699142937
transform -1 0 8832 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_227
timestamp 1699142937
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 1699142937
transform -1 0 8832 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_228
timestamp 1699142937
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 1699142937
transform -1 0 8832 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_229
timestamp 1699142937
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 1699142937
transform -1 0 8832 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_230
timestamp 1699142937
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 1699142937
transform -1 0 8832 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_231
timestamp 1699142937
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 1699142937
transform -1 0 8832 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_232
timestamp 1699142937
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 1699142937
transform -1 0 8832 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_233
timestamp 1699142937
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 1699142937
transform -1 0 8832 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_234
timestamp 1699142937
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 1699142937
transform -1 0 8832 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_235
timestamp 1699142937
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 1699142937
transform -1 0 8832 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_236
timestamp 1699142937
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 1699142937
transform -1 0 8832 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_237
timestamp 1699142937
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 1699142937
transform -1 0 8832 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_238
timestamp 1699142937
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 1699142937
transform -1 0 8832 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_239
timestamp 1699142937
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 1699142937
transform -1 0 8832 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_240
timestamp 1699142937
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 1699142937
transform -1 0 8832 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Left_241
timestamp 1699142937
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Right_102
timestamp 1699142937
transform -1 0 8832 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Left_242
timestamp 1699142937
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Right_103
timestamp 1699142937
transform -1 0 8832 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Left_243
timestamp 1699142937
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Right_104
timestamp 1699142937
transform -1 0 8832 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Left_244
timestamp 1699142937
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Right_105
timestamp 1699142937
transform -1 0 8832 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Left_245
timestamp 1699142937
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Right_106
timestamp 1699142937
transform -1 0 8832 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Left_246
timestamp 1699142937
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Right_107
timestamp 1699142937
transform -1 0 8832 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Left_247
timestamp 1699142937
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Right_108
timestamp 1699142937
transform -1 0 8832 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Left_248
timestamp 1699142937
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Right_109
timestamp 1699142937
transform -1 0 8832 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Left_249
timestamp 1699142937
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Right_110
timestamp 1699142937
transform -1 0 8832 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Left_250
timestamp 1699142937
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Right_111
timestamp 1699142937
transform -1 0 8832 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Left_251
timestamp 1699142937
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Right_112
timestamp 1699142937
transform -1 0 8832 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Left_252
timestamp 1699142937
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Right_113
timestamp 1699142937
transform -1 0 8832 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Left_253
timestamp 1699142937
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Right_114
timestamp 1699142937
transform -1 0 8832 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Left_254
timestamp 1699142937
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Right_115
timestamp 1699142937
transform -1 0 8832 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Left_255
timestamp 1699142937
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Right_116
timestamp 1699142937
transform -1 0 8832 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_256
timestamp 1699142937
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_117
timestamp 1699142937
transform -1 0 8832 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_257
timestamp 1699142937
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_118
timestamp 1699142937
transform -1 0 8832 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_258
timestamp 1699142937
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_119
timestamp 1699142937
transform -1 0 8832 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_259
timestamp 1699142937
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_120
timestamp 1699142937
transform -1 0 8832 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_260
timestamp 1699142937
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_121
timestamp 1699142937
transform -1 0 8832 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_261
timestamp 1699142937
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_122
timestamp 1699142937
transform -1 0 8832 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_262
timestamp 1699142937
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_123
timestamp 1699142937
transform -1 0 8832 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_263
timestamp 1699142937
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_124
timestamp 1699142937
transform -1 0 8832 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_264
timestamp 1699142937
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_125
timestamp 1699142937
transform -1 0 8832 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_265
timestamp 1699142937
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_126
timestamp 1699142937
transform -1 0 8832 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_266
timestamp 1699142937
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_127
timestamp 1699142937
transform -1 0 8832 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Left_267
timestamp 1699142937
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Right_128
timestamp 1699142937
transform -1 0 8832 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Left_268
timestamp 1699142937
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Right_129
timestamp 1699142937
transform -1 0 8832 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Left_269
timestamp 1699142937
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Right_130
timestamp 1699142937
transform -1 0 8832 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Left_270
timestamp 1699142937
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Right_131
timestamp 1699142937
transform -1 0 8832 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Left_271
timestamp 1699142937
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Right_132
timestamp 1699142937
transform -1 0 8832 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Left_272
timestamp 1699142937
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Right_133
timestamp 1699142937
transform -1 0 8832 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Left_273
timestamp 1699142937
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Right_134
timestamp 1699142937
transform -1 0 8832 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Left_274
timestamp 1699142937
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Right_135
timestamp 1699142937
transform -1 0 8832 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Left_275
timestamp 1699142937
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Right_136
timestamp 1699142937
transform -1 0 8832 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Left_276
timestamp 1699142937
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Right_137
timestamp 1699142937
transform -1 0 8832 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Left_277
timestamp 1699142937
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Right_138
timestamp 1699142937
transform -1 0 8832 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_278
timestamp 1699142937
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_279
timestamp 1699142937
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_280
timestamp 1699142937
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_281
timestamp 1699142937
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_282
timestamp 1699142937
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_283
timestamp 1699142937
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_284
timestamp 1699142937
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_285
timestamp 1699142937
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_286
timestamp 1699142937
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_287
timestamp 1699142937
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_288
timestamp 1699142937
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_289
timestamp 1699142937
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_290
timestamp 1699142937
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_291
timestamp 1699142937
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_292
timestamp 1699142937
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_293
timestamp 1699142937
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_294
timestamp 1699142937
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_295
timestamp 1699142937
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_296
timestamp 1699142937
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_297
timestamp 1699142937
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_298
timestamp 1699142937
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_299
timestamp 1699142937
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_300
timestamp 1699142937
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_301
timestamp 1699142937
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_302
timestamp 1699142937
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_303
timestamp 1699142937
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_304
timestamp 1699142937
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_305
timestamp 1699142937
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_306
timestamp 1699142937
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_307
timestamp 1699142937
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_308
timestamp 1699142937
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_309
timestamp 1699142937
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_310
timestamp 1699142937
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_311
timestamp 1699142937
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_312
timestamp 1699142937
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_313
timestamp 1699142937
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_314
timestamp 1699142937
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_315
timestamp 1699142937
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_316
timestamp 1699142937
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_317
timestamp 1699142937
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_318
timestamp 1699142937
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_319
timestamp 1699142937
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_320
timestamp 1699142937
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_321
timestamp 1699142937
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_322
timestamp 1699142937
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp 1699142937
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_324
timestamp 1699142937
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_325
timestamp 1699142937
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_326
timestamp 1699142937
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_327
timestamp 1699142937
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_328
timestamp 1699142937
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_329
timestamp 1699142937
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_330
timestamp 1699142937
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_331
timestamp 1699142937
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_332
timestamp 1699142937
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_333
timestamp 1699142937
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_334
timestamp 1699142937
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_335
timestamp 1699142937
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_336
timestamp 1699142937
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_337
timestamp 1699142937
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_338
timestamp 1699142937
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_339
timestamp 1699142937
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_340
timestamp 1699142937
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_341
timestamp 1699142937
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_342
timestamp 1699142937
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_343
timestamp 1699142937
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_344
timestamp 1699142937
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_345
timestamp 1699142937
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_346
timestamp 1699142937
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_347
timestamp 1699142937
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_348
timestamp 1699142937
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_349
timestamp 1699142937
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_350
timestamp 1699142937
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_351
timestamp 1699142937
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_352
timestamp 1699142937
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_353
timestamp 1699142937
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_354
timestamp 1699142937
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_355
timestamp 1699142937
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_356
timestamp 1699142937
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_357
timestamp 1699142937
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_358
timestamp 1699142937
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_359
timestamp 1699142937
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_360
timestamp 1699142937
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_361
timestamp 1699142937
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_362
timestamp 1699142937
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_363
timestamp 1699142937
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_364
timestamp 1699142937
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_365
timestamp 1699142937
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_366
timestamp 1699142937
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_367
timestamp 1699142937
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_368
timestamp 1699142937
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_369
timestamp 1699142937
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_370
timestamp 1699142937
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_371
timestamp 1699142937
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_372
timestamp 1699142937
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_373
timestamp 1699142937
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_374
timestamp 1699142937
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_375
timestamp 1699142937
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_376
timestamp 1699142937
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_377
timestamp 1699142937
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_378
timestamp 1699142937
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_379
timestamp 1699142937
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_380
timestamp 1699142937
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_381
timestamp 1699142937
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_382
timestamp 1699142937
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_383
timestamp 1699142937
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_384
timestamp 1699142937
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_385
timestamp 1699142937
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_386
timestamp 1699142937
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_387
timestamp 1699142937
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_388
timestamp 1699142937
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_389
timestamp 1699142937
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_390
timestamp 1699142937
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_391
timestamp 1699142937
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_392
timestamp 1699142937
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_393
timestamp 1699142937
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_394
timestamp 1699142937
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_395
timestamp 1699142937
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_396
timestamp 1699142937
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_397
timestamp 1699142937
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_398
timestamp 1699142937
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_399
timestamp 1699142937
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_400
timestamp 1699142937
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_401
timestamp 1699142937
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_402
timestamp 1699142937
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_403
timestamp 1699142937
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_404
timestamp 1699142937
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_405
timestamp 1699142937
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_406
timestamp 1699142937
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_407
timestamp 1699142937
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_408
timestamp 1699142937
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_409
timestamp 1699142937
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_410
timestamp 1699142937
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_411
timestamp 1699142937
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_412
timestamp 1699142937
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_413
timestamp 1699142937
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_414
timestamp 1699142937
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_415
timestamp 1699142937
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_416
timestamp 1699142937
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_417
timestamp 1699142937
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_418
timestamp 1699142937
transform 1 0 6256 0 1 77248
box -38 -48 130 592
<< labels >>
rlabel metal1 s 4968 77792 4968 77792 4 VDD
rlabel metal1 s 4968 77248 4968 77248 4 VSS
rlabel metal1 s 3992 6970 3992 6970 4 _000_
rlabel metal1 s 6762 16626 6762 16626 4 _001_
rlabel metal1 s 6854 18360 6854 18360 4 _002_
rlabel metal1 s 6808 19414 6808 19414 4 _003_
rlabel metal1 s 7176 20570 7176 20570 4 _004_
rlabel metal1 s 7912 21930 7912 21930 4 _005_
rlabel metal1 s 6808 23018 6808 23018 4 _006_
rlabel metal1 s 6762 24718 6762 24718 4 _007_
rlabel metal1 s 8142 25976 8142 25976 4 _008_
rlabel metal1 s 6302 26010 6302 26010 4 _009_
rlabel metal1 s 4370 7446 4370 7446 4 _010_
rlabel metal1 s 5842 7514 5842 7514 4 _011_
rlabel metal1 s 6762 7310 6762 7310 4 _012_
rlabel metal2 s 6854 8602 6854 8602 4 _013_
rlabel metal1 s 7038 10098 7038 10098 4 _014_
rlabel metal2 s 6854 11356 6854 11356 4 _015_
rlabel metal1 s 6808 12886 6808 12886 4 _016_
rlabel metal1 s 6900 13974 6900 13974 4 _017_
rlabel metal1 s 8004 15538 8004 15538 4 _018_
rlabel metal1 s 5152 42330 5152 42330 4 _019_
rlabel metal2 s 7038 33490 7038 33490 4 _020_
rlabel metal1 s 6785 34918 6785 34918 4 _021_
rlabel metal1 s 6785 36890 6785 36890 4 _022_
rlabel metal1 s 6785 37978 6785 37978 4 _023_
rlabel metal1 s 7636 39066 7636 39066 4 _024_
rlabel metal2 s 6946 40664 6946 40664 4 _025_
rlabel metal1 s 7360 28186 7360 28186 4 _026_
rlabel metal1 s 6854 29546 6854 29546 4 _027_
rlabel metal1 s 6854 31382 6854 31382 4 _028_
rlabel metal1 s 6785 32538 6785 32538 4 _029_
rlabel metal1 s 6946 66062 6946 66062 4 _030_
rlabel metal1 s 7130 67354 7130 67354 4 _031_
rlabel metal1 s 6854 68714 6854 68714 4 _032_
rlabel metal2 s 7038 70686 7038 70686 4 _033_
rlabel metal1 s 7084 72114 7084 72114 4 _034_
rlabel metal1 s 7406 73338 7406 73338 4 _035_
rlabel metal1 s 7130 44506 7130 44506 4 _036_
rlabel metal1 s 6854 45866 6854 45866 4 _037_
rlabel metal1 s 6854 47702 6854 47702 4 _038_
rlabel metal1 s 7038 48824 7038 48824 4 _039_
rlabel metal1 s 6854 50354 6854 50354 4 _040_
rlabel metal1 s 7038 51272 7038 51272 4 _041_
rlabel metal1 s 6854 53006 6854 53006 4 _042_
rlabel metal1 s 6854 54094 6854 54094 4 _043_
rlabel metal1 s 7038 55624 7038 55624 4 _044_
rlabel metal2 s 7038 57052 7038 57052 4 _045_
rlabel metal1 s 6946 58446 6946 58446 4 _046_
rlabel metal1 s 6854 59670 6854 59670 4 _047_
rlabel metal2 s 7038 60894 7038 60894 4 _048_
rlabel metal1 s 7038 62152 7038 62152 4 _049_
rlabel metal1 s 6716 64022 6716 64022 4 _050_
rlabel metal2 s 7038 64668 7038 64668 4 _051_
rlabel metal1 s 6893 42874 6893 42874 4 _052_
rlabel metal1 s 5375 34170 5375 34170 4 _053_
rlabel metal1 s 4968 35122 4968 35122 4 _054_
rlabel metal1 s 4922 36822 4922 36822 4 _055_
rlabel metal1 s 5014 37978 5014 37978 4 _056_
rlabel metal1 s 5106 39066 5106 39066 4 _057_
rlabel metal2 s 4738 28458 4738 28458 4 _058_
rlabel metal1 s 5152 28594 5152 28594 4 _059_
rlabel metal1 s 5152 30362 5152 30362 4 _060_
rlabel metal1 s 4922 31994 4922 31994 4 _061_
rlabel metal1 s 5382 65178 5382 65178 4 _062_
rlabel metal1 s 5198 66266 5198 66266 4 _063_
rlabel metal1 s 5152 67762 5152 67762 4 _064_
rlabel metal1 s 4968 68986 4968 68986 4 _065_
rlabel metal1 s 4876 70550 4876 70550 4 _066_
rlabel metal1 s 5198 71706 5198 71706 4 _067_
rlabel metal1 s 5428 72794 5428 72794 4 _068_
rlabel metal1 s 4968 45050 4968 45050 4 _069_
rlabel metal1 s 4968 46138 4968 46138 4 _070_
rlabel metal1 s 4738 47736 4738 47736 4 _071_
rlabel metal1 s 5060 48858 5060 48858 4 _072_
rlabel metal1 s 4876 50354 4876 50354 4 _073_
rlabel metal1 s 4830 51578 4830 51578 4 _074_
rlabel metal1 s 4738 53176 4738 53176 4 _075_
rlabel metal1 s 4922 54298 4922 54298 4 _076_
rlabel metal1 s 4876 55794 4876 55794 4 _077_
rlabel metal1 s 4784 57018 4784 57018 4 _078_
rlabel metal1 s 4876 58106 4876 58106 4 _079_
rlabel metal1 s 4738 59704 4738 59704 4 _080_
rlabel metal1 s 4784 60826 4784 60826 4 _081_
rlabel metal1 s 4692 62322 4692 62322 4 _082_
rlabel metal1 s 4731 63546 4731 63546 4 _083_
rlabel metal2 s 5198 43996 5198 43996 4 _084_
rlabel metal1 s 4692 40698 4692 40698 4 _085_
rlabel metal1 s 8556 41582 8556 41582 4 _086_
rlabel metal1 s 3726 7412 3726 7412 4 _087_
rlabel metal1 s 5796 6970 5796 6970 4 _088_
rlabel metal1 s 7360 6970 7360 6970 4 _089_
rlabel metal1 s 6394 7446 6394 7446 4 _090_
rlabel metal1 s 7038 8976 7038 8976 4 _091_
rlabel metal1 s 7590 10642 7590 10642 4 _092_
rlabel metal1 s 7406 11730 7406 11730 4 _093_
rlabel metal1 s 6946 13362 6946 13362 4 _094_
rlabel metal1 s 7452 14382 7452 14382 4 _095_
rlabel metal1 s 7498 16082 7498 16082 4 _096_
rlabel metal1 s 7406 17170 7406 17170 4 _097_
rlabel metal1 s 7590 18734 7590 18734 4 _098_
rlabel metal1 s 7038 19856 7038 19856 4 _099_
rlabel metal1 s 7406 20468 7406 20468 4 _100_
rlabel metal1 s 7222 22678 7222 22678 4 _101_
rlabel metal1 s 6486 23732 6486 23732 4 _102_
rlabel metal1 s 6946 25194 6946 25194 4 _103_
rlabel metal1 s 8280 26962 8280 26962 4 _104_
rlabel metal1 s 6394 25874 6394 25874 4 _105_
rlabel metal1 s 5566 42194 5566 42194 4 _106_
rlabel metal1 s 7360 45458 7360 45458 4 _107_
rlabel metal1 s 7590 39950 7590 39950 4 _108_
rlabel metal2 s 7222 33082 7222 33082 4 _109_
rlabel metal1 s 6624 33626 6624 33626 4 _110_
rlabel metal1 s 6578 36346 6578 36346 4 _111_
rlabel metal1 s 6624 37434 6624 37434 4 _112_
rlabel metal1 s 7636 38930 7636 38930 4 _113_
rlabel metal1 s 6624 40154 6624 40154 4 _114_
rlabel metal1 s 7728 28050 7728 28050 4 _115_
rlabel metal1 s 6670 29274 6670 29274 4 _116_
rlabel metal1 s 6624 30906 6624 30906 4 _117_
rlabel metal1 s 6624 31994 6624 31994 4 _118_
rlabel metal3 s 7383 60588 7383 60588 4 _119_
rlabel metal1 s 6486 66164 6486 66164 4 _120_
rlabel metal1 s 7590 67218 7590 67218 4 _121_
rlabel metal1 s 6578 68782 6578 68782 4 _122_
rlabel metal1 s 7084 70958 7084 70958 4 _123_
rlabel metal1 s 7130 71706 7130 71706 4 _124_
rlabel metal1 s 7728 73134 7728 73134 4 _125_
rlabel metal1 s 7084 44370 7084 44370 4 _126_
rlabel metal1 s 6486 45968 6486 45968 4 _127_
rlabel metal1 s 6670 47226 6670 47226 4 _128_
rlabel metal1 s 7682 48314 7682 48314 4 _129_
rlabel metal1 s 7222 52564 7222 52564 4 _130_
rlabel metal1 s 6578 49402 6578 49402 4 _131_
rlabel metal1 s 6578 51034 6578 51034 4 _132_
rlabel metal1 s 6578 52666 6578 52666 4 _133_
rlabel metal1 s 6578 53754 6578 53754 4 _134_
rlabel metal1 s 6578 55386 6578 55386 4 _135_
rlabel metal1 s 6808 56474 6808 56474 4 _136_
rlabel metal1 s 6624 58106 6624 58106 4 _137_
rlabel metal1 s 6624 59194 6624 59194 4 _138_
rlabel metal1 s 6762 60282 6762 60282 4 _139_
rlabel metal1 s 6624 61914 6624 61914 4 _140_
rlabel metal1 s 6440 63546 6440 63546 4 _141_
rlabel metal1 s 7176 63478 7176 63478 4 _142_
rlabel metal1 s 7268 42330 7268 42330 4 _143_
rlabel metal2 s 5474 34102 5474 34102 4 _144_
rlabel metal1 s 5382 35666 5382 35666 4 _145_
rlabel metal1 s 5336 37230 5336 37230 4 _146_
rlabel metal1 s 5382 37842 5382 37842 4 _147_
rlabel metal1 s 5428 38930 5428 38930 4 _148_
rlabel metal1 s 5198 29138 5198 29138 4 _149_
rlabel metal1 s 5428 29138 5428 29138 4 _150_
rlabel metal1 s 5888 30226 5888 30226 4 _151_
rlabel metal1 s 5428 31790 5428 31790 4 _152_
rlabel metal1 s 5842 65076 5842 65076 4 _153_
rlabel metal1 s 5934 66130 5934 66130 4 _154_
rlabel metal1 s 5428 68306 5428 68306 4 _155_
rlabel metal1 s 5474 68782 5474 68782 4 _156_
rlabel metal1 s 5474 70958 5474 70958 4 _157_
rlabel metal1 s 5934 71570 5934 71570 4 _158_
rlabel metal1 s 6026 72658 6026 72658 4 _159_
rlabel metal1 s 5566 44846 5566 44846 4 _160_
rlabel metal1 s 5428 45934 5428 45934 4 _161_
rlabel metal1 s 5428 48110 5428 48110 4 _162_
rlabel metal1 s 5382 48722 5382 48722 4 _163_
rlabel metal1 s 5290 50898 5290 50898 4 _164_
rlabel metal1 s 5198 51374 5198 51374 4 _165_
rlabel metal1 s 5244 53550 5244 53550 4 _166_
rlabel metal1 s 5244 54162 5244 54162 4 _167_
rlabel metal1 s 5244 56338 5244 56338 4 _168_
rlabel metal1 s 5060 56814 5060 56814 4 _169_
rlabel metal1 s 5244 57902 5244 57902 4 _170_
rlabel metal1 s 5152 60078 5152 60078 4 _171_
rlabel metal1 s 5106 60554 5106 60554 4 _172_
rlabel metal1 s 5106 62866 5106 62866 4 _173_
rlabel metal1 s 5152 63954 5152 63954 4 _174_
rlabel metal2 s 5382 43894 5382 43894 4 _175_
rlabel metal1 s 5060 40154 5060 40154 4 _176_
rlabel metal1 s 7682 33082 7682 33082 4 adc_cfg1[0]
rlabel metal2 s 8418 66725 8418 66725 4 adc_cfg1[10]
rlabel metal2 s 8418 67949 8418 67949 4 adc_cfg1[11]
rlabel metal3 s 8418 69173 8418 69173 4 adc_cfg1[12]
rlabel metal2 s 8418 70669 8418 70669 4 adc_cfg1[13]
rlabel metal1 s 8464 71706 8464 71706 4 adc_cfg1[14]
rlabel metal2 s 8418 73661 8418 73661 4 adc_cfg1[15]
rlabel metal2 s 8418 35309 8418 35309 4 adc_cfg1[1]
rlabel metal2 s 8418 36431 8418 36431 4 adc_cfg1[2]
rlabel metal2 s 8418 38029 8418 38029 4 adc_cfg1[3]
rlabel metal2 s 8418 39151 8418 39151 4 adc_cfg1[4]
rlabel metal2 s 8418 40749 8418 40749 4 adc_cfg1[5]
rlabel metal2 s 8418 28271 8418 28271 4 adc_cfg1[6]
rlabel metal2 s 8418 29869 8418 29869 4 adc_cfg1[7]
rlabel metal2 s 8418 30991 8418 30991 4 adc_cfg1[8]
rlabel metal1 s 8464 32742 8464 32742 4 adc_cfg1[9]
rlabel metal2 s 8418 44591 8418 44591 4 adc_cfg2[0]
rlabel metal1 s 8464 58854 8464 58854 4 adc_cfg2[10]
rlabel metal2 s 8418 59789 8418 59789 4 adc_cfg2[11]
rlabel metal3 s 8418 61013 8418 61013 4 adc_cfg2[12]
rlabel metal2 s 8418 62509 8418 62509 4 adc_cfg2[13]
rlabel metal1 s 8418 63512 8418 63512 4 adc_cfg2[14]
rlabel metal2 s 8418 65229 8418 65229 4 adc_cfg2[15]
rlabel metal2 s 8418 46189 8418 46189 4 adc_cfg2[1]
rlabel metal2 s 8418 47311 8418 47311 4 adc_cfg2[2]
rlabel metal2 s 8418 48909 8418 48909 4 adc_cfg2[3]
rlabel metal2 s 8418 50031 8418 50031 4 adc_cfg2[4]
rlabel metal2 s 8418 51629 8418 51629 4 adc_cfg2[5]
rlabel metal2 s 8418 52751 8418 52751 4 adc_cfg2[6]
rlabel metal2 s 8418 54349 8418 54349 4 adc_cfg2[7]
rlabel metal1 s 7912 54842 7912 54842 4 adc_cfg2[8]
rlabel metal1 s 8326 57222 8326 57222 4 adc_cfg2[9]
rlabel metal2 s 6578 33694 6578 33694 4 adc_cfg_load_r\[0\]
rlabel metal1 s 6762 66810 6762 66810 4 adc_cfg_load_r\[10\]
rlabel metal2 s 6578 68102 6578 68102 4 adc_cfg_load_r\[11\]
rlabel metal1 s 6762 69326 6762 69326 4 adc_cfg_load_r\[12\]
rlabel metal1 s 6118 70822 6118 70822 4 adc_cfg_load_r\[13\]
rlabel metal1 s 6394 71502 6394 71502 4 adc_cfg_load_r\[14\]
rlabel metal2 s 6854 72148 6854 72148 4 adc_cfg_load_r\[15\]
rlabel metal1 s 6716 72658 6716 72658 4 adc_cfg_load_r\[16\]
rlabel metal1 s 6762 46478 6762 46478 4 adc_cfg_load_r\[17\]
rlabel metal1 s 5980 47022 5980 47022 4 adc_cfg_load_r\[18\]
rlabel metal1 s 6486 48110 6486 48110 4 adc_cfg_load_r\[19\]
rlabel metal1 s 6164 35258 6164 35258 4 adc_cfg_load_r\[1\]
rlabel metal1 s 6072 50490 6072 50490 4 adc_cfg_load_r\[20\]
rlabel metal2 s 5750 51612 5750 51612 4 adc_cfg_load_r\[21\]
rlabel metal2 s 6210 52122 6210 52122 4 adc_cfg_load_r\[22\]
rlabel metal1 s 6394 53482 6394 53482 4 adc_cfg_load_r\[23\]
rlabel metal1 s 5980 55590 5980 55590 4 adc_cfg_load_r\[24\]
rlabel metal1 s 6440 56406 6440 56406 4 adc_cfg_load_r\[25\]
rlabel metal1 s 6118 58310 6118 58310 4 adc_cfg_load_r\[26\]
rlabel metal2 s 6210 59228 6210 59228 4 adc_cfg_load_r\[27\]
rlabel metal1 s 6348 60010 6348 60010 4 adc_cfg_load_r\[28\]
rlabel metal2 s 6118 61472 6118 61472 4 adc_cfg_load_r\[29\]
rlabel metal2 s 6210 36992 6210 36992 4 adc_cfg_load_r\[2\]
rlabel metal1 s 5934 63546 5934 63546 4 adc_cfg_load_r\[30\]
rlabel metal1 s 6486 55250 6486 55250 4 adc_cfg_load_r\[31\]
rlabel metal1 s 6164 41242 6164 41242 4 adc_cfg_load_r\[32\]
rlabel metal2 s 5934 37468 5934 37468 4 adc_cfg_load_r\[3\]
rlabel metal2 s 5934 38454 5934 38454 4 adc_cfg_load_r\[4\]
rlabel metal1 s 6072 38998 6072 38998 4 adc_cfg_load_r\[5\]
rlabel metal2 s 6578 28254 6578 28254 4 adc_cfg_load_r\[6\]
rlabel metal1 s 6578 29206 6578 29206 4 adc_cfg_load_r\[7\]
rlabel metal1 s 6118 31654 6118 31654 4 adc_cfg_load_r\[8\]
rlabel metal2 s 7130 40324 7130 40324 4 adc_cfg_load_r\[9\]
rlabel metal1 s 6808 42534 6808 42534 4 adc_cfg_written_r
rlabel metal1 s 7498 42126 7498 42126 4 adc_conv_finished
rlabel metal1 s 8694 43758 8694 43758 4 adc_conv_finished_osr
rlabel metal1 s 8694 5678 8694 5678 4 adc_res[0]
rlabel metal1 s 6578 19788 6578 19788 4 adc_res[10]
rlabel metal1 s 6762 21556 6762 21556 4 adc_res[11]
rlabel metal1 s 6946 22576 6946 22576 4 adc_res[12]
rlabel metal1 s 7406 22610 7406 22610 4 adc_res[13]
rlabel metal1 s 8096 27438 8096 27438 4 adc_res[14]
rlabel metal1 s 8694 27438 8694 27438 4 adc_res[15]
rlabel metal1 s 7268 9554 7268 9554 4 adc_res[1]
rlabel metal1 s 6578 8908 6578 8908 4 adc_res[2]
rlabel metal1 s 7728 12206 7728 12206 4 adc_res[3]
rlabel metal1 s 6578 11662 6578 11662 4 adc_res[4]
rlabel metal1 s 6486 13260 6486 13260 4 adc_res[5]
rlabel metal1 s 8694 14994 8694 14994 4 adc_res[6]
rlabel metal1 s 6670 17170 6670 17170 4 adc_res[7]
rlabel metal1 s 7820 17646 7820 17646 4 adc_res[8]
rlabel metal1 s 7728 20434 7728 20434 4 adc_res[9]
rlabel metal2 s 8326 16932 8326 16932 4 adc_res_r\[10\]
rlabel metal2 s 8418 17612 8418 17612 4 adc_res_r\[11\]
rlabel metal1 s 8602 19482 8602 19482 4 adc_res_r\[12\]
rlabel metal2 s 8418 20332 8418 20332 4 adc_res_r\[13\]
rlabel metal2 s 7038 21692 7038 21692 4 adc_res_r\[14\]
rlabel metal2 s 8326 23460 8326 23460 4 adc_res_r\[15\]
rlabel metal1 s 8418 23766 8418 23766 4 adc_res_r\[16\]
rlabel metal1 s 6854 25330 6854 25330 4 adc_res_r\[17\]
rlabel metal1 s 8004 26418 8004 26418 4 adc_res_r\[18\]
rlabel metal1 s 6394 26554 6394 26554 4 adc_res_r\[19\]
rlabel metal1 s 5888 7310 5888 7310 4 adc_res_r\[1\]
rlabel metal1 s 7268 7922 7268 7922 4 adc_res_r\[2\]
rlabel metal2 s 8418 6732 8418 6732 4 adc_res_r\[3\]
rlabel metal1 s 7774 8602 7774 8602 4 adc_res_r\[4\]
rlabel metal2 s 8418 9452 8418 9452 4 adc_res_r\[5\]
rlabel metal1 s 7774 11322 7774 11322 4 adc_res_r\[6\]
rlabel metal2 s 8326 12517 8326 12517 4 adc_res_r\[7\]
rlabel metal1 s 7498 13362 7498 13362 4 adc_res_r\[8\]
rlabel metal2 s 6670 15164 6670 15164 4 adc_res_r\[9\]
rlabel metal1 s 6670 40528 6670 40528 4 clk
rlabel metal1 s 6118 40358 6118 40358 4 clknet_0_clk
rlabel metal1 s 4554 38318 4554 38318 4 clknet_3_0_0_clk
rlabel metal2 s 6762 37230 6762 37230 4 clknet_3_1_0_clk
rlabel metal1 s 6348 12818 6348 12818 4 clknet_3_2_0_clk
rlabel metal1 s 7452 22066 7452 22066 4 clknet_3_3_0_clk
rlabel metal2 s 4462 52462 4462 52462 4 clknet_3_4_0_clk
rlabel metal1 s 4968 72114 4968 72114 4 clknet_3_5_0_clk
rlabel metal1 s 6440 56882 6440 56882 4 clknet_3_6_0_clk
rlabel metal1 s 5612 58446 5612 58446 4 clknet_3_7_0_clk
rlabel metal2 s 9154 1554 9154 1554 4 conv_finish
rlabel metal1 s 7866 42194 7866 42194 4 conv_finish_sel
rlabel metal2 s 5842 1588 5842 1588 4 dat_i
rlabel metal2 s 4186 1520 4186 1520 4 dat_o
rlabel metal2 s 7498 959 7498 959 4 load
rlabel metal1 s 7866 42330 7866 42330 4 net1
rlabel metal1 s 8050 7922 8050 7922 4 net10
rlabel metal2 s 6762 9316 6762 9316 4 net11
rlabel metal1 s 8004 10574 8004 10574 4 net12
rlabel metal2 s 6762 12002 6762 12002 4 net13
rlabel metal1 s 8234 13430 8234 13430 4 net14
rlabel metal2 s 8234 14620 8234 14620 4 net15
rlabel metal1 s 7590 16014 7590 16014 4 net16
rlabel metal1 s 7774 17714 7774 17714 4 net17
rlabel metal1 s 8004 18802 8004 18802 4 net18
rlabel metal4 s 6693 2652 6693 2652 4 net19
rlabel metal1 s 8050 42262 8050 42262 4 net2
rlabel metal1 s 7682 2618 7682 2618 4 net20
rlabel metal1 s 6394 40086 6394 40086 4 net21
rlabel metal2 s 7958 33728 7958 33728 4 net22
rlabel metal1 s 8280 66538 8280 66538 4 net23
rlabel metal1 s 7728 68306 7728 68306 4 net24
rlabel metal1 s 7728 69394 7728 69394 4 net25
rlabel metal1 s 8280 70414 8280 70414 4 net26
rlabel metal1 s 8050 71638 8050 71638 4 net27
rlabel metal1 s 8280 73542 8280 73542 4 net28
rlabel metal1 s 7820 34918 7820 34918 4 net29
rlabel metal1 s 8418 5882 8418 5882 4 net3
rlabel metal1 s 8556 36142 8556 36142 4 net30
rlabel metal1 s 7820 37638 7820 37638 4 net31
rlabel metal1 s 8556 38930 8556 38930 4 net32
rlabel metal1 s 8694 40358 8694 40358 4 net33
rlabel metal1 s 8556 28050 8556 28050 4 net34
rlabel metal1 s 8694 29478 8694 29478 4 net35
rlabel metal1 s 8556 30702 8556 30702 4 net36
rlabel metal1 s 7820 32198 7820 32198 4 net37
rlabel metal1 s 8694 45050 8694 45050 4 net38
rlabel metal1 s 7820 58310 7820 58310 4 net39
rlabel metal1 s 6992 19686 6992 19686 4 net4
rlabel metal1 s 7820 59398 7820 59398 4 net40
rlabel metal2 s 7774 60486 7774 60486 4 net41
rlabel metal1 s 7820 62118 7820 62118 4 net42
rlabel metal1 s 8188 63342 8188 63342 4 net43
rlabel metal1 s 8234 64294 8234 64294 4 net44
rlabel metal1 s 7728 46546 7728 46546 4 net45
rlabel metal1 s 8556 47022 8556 47022 4 net46
rlabel metal1 s 8280 48518 8280 48518 4 net47
rlabel metal1 s 8234 49776 8234 49776 4 net48
rlabel metal1 s 8234 51238 8234 51238 4 net49
rlabel metal1 s 7590 21658 7590 21658 4 net5
rlabel metal2 s 8234 52666 8234 52666 4 net50
rlabel metal1 s 7774 53958 7774 53958 4 net51
rlabel metal2 s 8510 55420 8510 55420 4 net52
rlabel metal1 s 7452 57426 7452 57426 4 net53
rlabel metal1 s 8050 2414 8050 2414 4 net54
rlabel metal1 s 5014 2414 5014 2414 4 net55
rlabel metal2 s 4830 7072 4830 7072 4 net56
rlabel metal2 s 7958 17731 7958 17731 4 net57
rlabel metal1 s 8004 30906 8004 30906 4 net58
rlabel metal1 s 6854 36652 6854 36652 4 net59
rlabel metal1 s 7820 22678 7820 22678 4 net6
rlabel metal1 s 6401 39338 6401 39338 4 net60
rlabel metal2 s 7130 40800 7130 40800 4 net61
rlabel metal1 s 8089 56814 8089 56814 4 net62
rlabel metal1 s 6532 56474 6532 56474 4 net63
rlabel metal1 s 5789 58514 5789 58514 4 net64
rlabel metal1 s 7307 70550 7307 70550 4 net65
rlabel metal1 s 6631 73066 6631 73066 4 net66
rlabel metal1 s 8418 13260 8418 13260 4 net67
rlabel metal1 s 8142 21454 8142 21454 4 net68
rlabel metal2 s 6118 34510 6118 34510 4 net69
rlabel metal1 s 7774 22474 7774 22474 4 net7
rlabel metal1 s 6072 37298 6072 37298 4 net70
rlabel metal2 s 6026 48909 6026 48909 4 net71
rlabel metal1 s 5888 60622 5888 60622 4 net72
rlabel metal1 s 6164 57018 6164 57018 4 net73
rlabel metal1 s 2392 3026 2392 3026 4 net74
rlabel metal2 s 1886 2754 1886 2754 4 net75
rlabel metal2 s 5106 8058 5106 8058 4 net76
rlabel metal1 s 6256 25738 6256 25738 4 net77
rlabel metal1 s 8004 22746 8004 22746 4 net78
rlabel metal1 s 8050 10778 8050 10778 4 net79
rlabel metal1 s 8050 25330 8050 25330 4 net8
rlabel metal1 s 8050 16218 8050 16218 4 net80
rlabel metal1 s 7912 13226 7912 13226 4 net81
rlabel metal1 s 7958 7854 7958 7854 4 net82
rlabel metal1 s 8004 18734 8004 18734 4 net83
rlabel metal1 s 8004 9146 8004 9146 4 net84
rlabel metal1 s 8004 20026 8004 20026 4 net85
rlabel metal2 s 7866 11968 7866 11968 4 net86
rlabel metal2 s 7866 17408 7866 17408 4 net87
rlabel metal1 s 8142 14484 8142 14484 4 net88
rlabel metal1 s 7912 21522 7912 21522 4 net89
rlabel metal1 s 8050 27030 8050 27030 4 net9
rlabel metal1 s 7912 25194 7912 25194 4 net90
rlabel metal2 s 7866 6528 7866 6528 4 net91
rlabel metal2 s 7774 26758 7774 26758 4 net92
rlabel metal1 s 6210 6868 6210 6868 4 net93
rlabel metal2 s 7866 23936 7866 23936 4 net94
rlabel metal1 s 7452 55250 7452 55250 4 net95
rlabel metal2 s 2714 77877 2714 77877 4 rst_n
rlabel metal2 s 2530 823 2530 823 4 tie0
rlabel metal2 s 874 1792 874 1792 4 tie1
flabel metal5 s -1076 73416 11012 73736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 68416 11012 68736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 63416 11012 63736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 58416 11012 58736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 53416 11012 53736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 48416 11012 48736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 43416 11012 43736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 38416 11012 38736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 33416 11012 33736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 28416 11012 28736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 23416 11012 23736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 18416 11012 18736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 13416 11012 13736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 8416 11012 8736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -1076 3416 11012 3736 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal4 s 7344 -4 7664 79972 0 FreeSans 2400 90 0 0 VDD
port 1 nsew
flabel metal4 s 2344 -4 2664 79972 0 FreeSans 2400 90 0 0 VDD
port 1 nsew
flabel metal4 s 10032 656 10352 79312 0 FreeSans 2400 90 0 0 VDD
port 1 nsew
flabel metal5 s -416 78992 10352 79312 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal5 s -416 656 10352 976 0 FreeSans 3200 0 0 0 VDD
port 1 nsew
flabel metal4 s -416 656 -96 79312 0 FreeSans 2400 90 0 0 VDD
port 1 nsew
flabel metal5 s -1076 74076 11012 74396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 69076 11012 69396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 64076 11012 64396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 59076 11012 59396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 54076 11012 54396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 49076 11012 49396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 44076 11012 44396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 39076 11012 39396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 34076 11012 34396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 29076 11012 29396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 24076 11012 24396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 19076 11012 19396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 14076 11012 14396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 9076 11012 9396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 4076 11012 4396 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal4 s 8004 -4 8324 79972 0 FreeSans 2400 90 0 0 VSS
port 2 nsew
flabel metal4 s 3004 -4 3324 79972 0 FreeSans 2400 90 0 0 VSS
port 2 nsew
flabel metal4 s 10692 -4 11012 79972 0 FreeSans 2400 90 0 0 VSS
port 2 nsew
flabel metal5 s -1076 79652 11012 79972 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal5 s -1076 -4 11012 316 0 FreeSans 3200 0 0 0 VSS
port 2 nsew
flabel metal4 s -1076 -4 -756 79972 0 FreeSans 2400 90 0 0 VSS
port 2 nsew
flabel metal3 s 9200 33736 10000 33856 0 FreeSans 600 0 0 0 adc_cfg1[0]
port 3 nsew
flabel metal3 s 9200 66376 10000 66496 0 FreeSans 600 0 0 0 adc_cfg1[10]
port 4 nsew
flabel metal3 s 9200 67736 10000 67856 0 FreeSans 600 0 0 0 adc_cfg1[11]
port 5 nsew
flabel metal3 s 9200 69096 10000 69216 0 FreeSans 600 0 0 0 adc_cfg1[12]
port 6 nsew
flabel metal3 s 9200 70456 10000 70576 0 FreeSans 600 0 0 0 adc_cfg1[13]
port 7 nsew
flabel metal3 s 9200 71816 10000 71936 0 FreeSans 600 0 0 0 adc_cfg1[14]
port 8 nsew
flabel metal3 s 9200 73176 10000 73296 0 FreeSans 600 0 0 0 adc_cfg1[15]
port 9 nsew
flabel metal3 s 9200 35096 10000 35216 0 FreeSans 600 0 0 0 adc_cfg1[1]
port 10 nsew
flabel metal3 s 9200 36456 10000 36576 0 FreeSans 600 0 0 0 adc_cfg1[2]
port 11 nsew
flabel metal3 s 9200 37816 10000 37936 0 FreeSans 600 0 0 0 adc_cfg1[3]
port 12 nsew
flabel metal3 s 9200 39176 10000 39296 0 FreeSans 600 0 0 0 adc_cfg1[4]
port 13 nsew
flabel metal3 s 9200 40536 10000 40656 0 FreeSans 600 0 0 0 adc_cfg1[5]
port 14 nsew
flabel metal3 s 9200 28296 10000 28416 0 FreeSans 600 0 0 0 adc_cfg1[6]
port 15 nsew
flabel metal3 s 9200 29656 10000 29776 0 FreeSans 600 0 0 0 adc_cfg1[7]
port 16 nsew
flabel metal3 s 9200 31016 10000 31136 0 FreeSans 600 0 0 0 adc_cfg1[8]
port 17 nsew
flabel metal3 s 9200 32376 10000 32496 0 FreeSans 600 0 0 0 adc_cfg1[9]
port 18 nsew
flabel metal3 s 9200 44616 10000 44736 0 FreeSans 600 0 0 0 adc_cfg2[0]
port 19 nsew
flabel metal3 s 9200 58216 10000 58336 0 FreeSans 600 0 0 0 adc_cfg2[10]
port 20 nsew
flabel metal3 s 9200 59576 10000 59696 0 FreeSans 600 0 0 0 adc_cfg2[11]
port 21 nsew
flabel metal3 s 9200 60936 10000 61056 0 FreeSans 600 0 0 0 adc_cfg2[12]
port 22 nsew
flabel metal3 s 9200 62296 10000 62416 0 FreeSans 600 0 0 0 adc_cfg2[13]
port 23 nsew
flabel metal3 s 9200 63656 10000 63776 0 FreeSans 600 0 0 0 adc_cfg2[14]
port 24 nsew
flabel metal3 s 9200 65016 10000 65136 0 FreeSans 600 0 0 0 adc_cfg2[15]
port 25 nsew
flabel metal3 s 9200 45976 10000 46096 0 FreeSans 600 0 0 0 adc_cfg2[1]
port 26 nsew
flabel metal3 s 9200 47336 10000 47456 0 FreeSans 600 0 0 0 adc_cfg2[2]
port 27 nsew
flabel metal3 s 9200 48696 10000 48816 0 FreeSans 600 0 0 0 adc_cfg2[3]
port 28 nsew
flabel metal3 s 9200 50056 10000 50176 0 FreeSans 600 0 0 0 adc_cfg2[4]
port 29 nsew
flabel metal3 s 9200 51416 10000 51536 0 FreeSans 600 0 0 0 adc_cfg2[5]
port 30 nsew
flabel metal3 s 9200 52776 10000 52896 0 FreeSans 600 0 0 0 adc_cfg2[6]
port 31 nsew
flabel metal3 s 9200 54136 10000 54256 0 FreeSans 600 0 0 0 adc_cfg2[7]
port 32 nsew
flabel metal3 s 9200 55496 10000 55616 0 FreeSans 600 0 0 0 adc_cfg2[8]
port 33 nsew
flabel metal3 s 9200 56856 10000 56976 0 FreeSans 600 0 0 0 adc_cfg2[9]
port 34 nsew
flabel metal3 s 9200 41896 10000 42016 0 FreeSans 600 0 0 0 adc_conv_finished
port 35 nsew
flabel metal3 s 9200 43256 10000 43376 0 FreeSans 600 0 0 0 adc_conv_finished_osr
port 36 nsew
flabel metal3 s 9200 6536 10000 6656 0 FreeSans 600 0 0 0 adc_res[0]
port 37 nsew
flabel metal3 s 9200 20136 10000 20256 0 FreeSans 600 0 0 0 adc_res[10]
port 38 nsew
flabel metal3 s 9200 21496 10000 21616 0 FreeSans 600 0 0 0 adc_res[11]
port 39 nsew
flabel metal3 s 9200 22856 10000 22976 0 FreeSans 600 0 0 0 adc_res[12]
port 40 nsew
flabel metal3 s 9200 24216 10000 24336 0 FreeSans 600 0 0 0 adc_res[13]
port 41 nsew
flabel metal3 s 9200 25576 10000 25696 0 FreeSans 600 0 0 0 adc_res[14]
port 42 nsew
flabel metal3 s 9200 26936 10000 27056 0 FreeSans 600 0 0 0 adc_res[15]
port 43 nsew
flabel metal3 s 9200 7896 10000 8016 0 FreeSans 600 0 0 0 adc_res[1]
port 44 nsew
flabel metal3 s 9200 9256 10000 9376 0 FreeSans 600 0 0 0 adc_res[2]
port 45 nsew
flabel metal3 s 9200 10616 10000 10736 0 FreeSans 600 0 0 0 adc_res[3]
port 46 nsew
flabel metal3 s 9200 11976 10000 12096 0 FreeSans 600 0 0 0 adc_res[4]
port 47 nsew
flabel metal3 s 9200 13336 10000 13456 0 FreeSans 600 0 0 0 adc_res[5]
port 48 nsew
flabel metal3 s 9200 14696 10000 14816 0 FreeSans 600 0 0 0 adc_res[6]
port 49 nsew
flabel metal3 s 9200 16056 10000 16176 0 FreeSans 600 0 0 0 adc_res[7]
port 50 nsew
flabel metal3 s 9200 17416 10000 17536 0 FreeSans 600 0 0 0 adc_res[8]
port 51 nsew
flabel metal3 s 9200 18776 10000 18896 0 FreeSans 600 0 0 0 adc_res[9]
port 52 nsew
flabel metal2 s 7470 79200 7526 80000 0 FreeSans 280 90 0 0 clk
port 53 nsew
flabel metal2 s 9126 0 9182 800 0 FreeSans 280 90 0 0 conv_finish
port 54 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 dat_i
port 55 nsew
flabel metal2 s 4158 0 4214 800 0 FreeSans 280 90 0 0 dat_o
port 56 nsew
flabel metal2 s 7470 0 7526 800 0 FreeSans 280 90 0 0 load
port 57 nsew
flabel metal2 s 2502 79200 2558 80000 0 FreeSans 280 90 0 0 rst_n
port 58 nsew
flabel metal2 s 2502 0 2558 800 0 FreeSans 280 90 0 0 tie0
port 59 nsew
flabel metal2 s 846 0 902 800 0 FreeSans 280 90 0 0 tie1
port 60 nsew
<< properties >>
string FIXED_BBOX 0 0 10000 80000
string GDS_END 1226772
string GDS_FILE adc_bridge.gds
string GDS_START 153194
<< end >>
