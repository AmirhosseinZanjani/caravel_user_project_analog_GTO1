magic
tech sky130A
timestamp 1694531879
use PA_nfet_w15_l015  PA_nfet_w15_l015_0
timestamp 1694529803
transform 1 0 902 0 1 123
box -61 -123 779 595
use PA_nfet_w15_l015  PA_nfet_w15_l015_1
timestamp 1694529803
transform 1 0 116 0 1 123
box -61 -123 779 595
<< end >>
