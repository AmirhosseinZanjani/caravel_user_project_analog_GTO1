magic
tech sky130A
magscale 1 2
timestamp 1692605656
<< error_p >>
rect -29 1020 29 1026
rect -29 986 -17 1020
rect -29 980 29 986
rect -29 826 29 832
rect -29 792 -17 826
rect -29 786 29 792
rect -29 718 29 724
rect -29 684 -17 718
rect -29 678 29 684
rect -29 524 29 530
rect -29 490 -17 524
rect -29 484 29 490
rect -29 416 29 422
rect -29 382 -17 416
rect -29 376 29 382
rect -29 222 29 228
rect -29 188 -17 222
rect -29 182 29 188
rect -29 114 29 120
rect -29 80 -17 114
rect -29 74 29 80
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect -29 -120 29 -114
rect -29 -188 29 -182
rect -29 -222 -17 -188
rect -29 -228 29 -222
rect -29 -382 29 -376
rect -29 -416 -17 -382
rect -29 -422 29 -416
rect -29 -490 29 -484
rect -29 -524 -17 -490
rect -29 -530 29 -524
rect -29 -684 29 -678
rect -29 -718 -17 -684
rect -29 -724 29 -718
rect -29 -792 29 -786
rect -29 -826 -17 -792
rect -29 -832 29 -826
rect -29 -986 29 -980
rect -29 -1020 -17 -986
rect -29 -1026 29 -1020
<< pwell >>
rect -211 -1158 211 1158
<< nmos >>
rect -15 864 15 948
rect -15 562 15 646
rect -15 260 15 344
rect -15 -42 15 42
rect -15 -344 15 -260
rect -15 -646 15 -562
rect -15 -948 15 -864
<< ndiff >>
rect -73 936 -15 948
rect -73 876 -61 936
rect -27 876 -15 936
rect -73 864 -15 876
rect 15 936 73 948
rect 15 876 27 936
rect 61 876 73 936
rect 15 864 73 876
rect -73 634 -15 646
rect -73 574 -61 634
rect -27 574 -15 634
rect -73 562 -15 574
rect 15 634 73 646
rect 15 574 27 634
rect 61 574 73 634
rect 15 562 73 574
rect -73 332 -15 344
rect -73 272 -61 332
rect -27 272 -15 332
rect -73 260 -15 272
rect 15 332 73 344
rect 15 272 27 332
rect 61 272 73 332
rect 15 260 73 272
rect -73 30 -15 42
rect -73 -30 -61 30
rect -27 -30 -15 30
rect -73 -42 -15 -30
rect 15 30 73 42
rect 15 -30 27 30
rect 61 -30 73 30
rect 15 -42 73 -30
rect -73 -272 -15 -260
rect -73 -332 -61 -272
rect -27 -332 -15 -272
rect -73 -344 -15 -332
rect 15 -272 73 -260
rect 15 -332 27 -272
rect 61 -332 73 -272
rect 15 -344 73 -332
rect -73 -574 -15 -562
rect -73 -634 -61 -574
rect -27 -634 -15 -574
rect -73 -646 -15 -634
rect 15 -574 73 -562
rect 15 -634 27 -574
rect 61 -634 73 -574
rect 15 -646 73 -634
rect -73 -876 -15 -864
rect -73 -936 -61 -876
rect -27 -936 -15 -876
rect -73 -948 -15 -936
rect 15 -876 73 -864
rect 15 -936 27 -876
rect 61 -936 73 -876
rect 15 -948 73 -936
<< ndiffc >>
rect -61 876 -27 936
rect 27 876 61 936
rect -61 574 -27 634
rect 27 574 61 634
rect -61 272 -27 332
rect 27 272 61 332
rect -61 -30 -27 30
rect 27 -30 61 30
rect -61 -332 -27 -272
rect 27 -332 61 -272
rect -61 -634 -27 -574
rect 27 -634 61 -574
rect -61 -936 -27 -876
rect 27 -936 61 -876
<< psubdiff >>
rect -175 1088 -79 1122
rect 79 1088 175 1122
rect -175 1026 -141 1088
rect 141 1026 175 1088
rect -175 -1088 -141 -1026
rect 141 -1088 175 -1026
rect -175 -1122 -79 -1088
rect 79 -1122 175 -1088
<< psubdiffcont >>
rect -79 1088 79 1122
rect -175 -1026 -141 1026
rect 141 -1026 175 1026
rect -79 -1122 79 -1088
<< poly >>
rect -33 1020 33 1036
rect -33 986 -17 1020
rect 17 986 33 1020
rect -33 970 33 986
rect -15 948 15 970
rect -15 842 15 864
rect -33 826 33 842
rect -33 792 -17 826
rect 17 792 33 826
rect -33 776 33 792
rect -33 718 33 734
rect -33 684 -17 718
rect 17 684 33 718
rect -33 668 33 684
rect -15 646 15 668
rect -15 540 15 562
rect -33 524 33 540
rect -33 490 -17 524
rect 17 490 33 524
rect -33 474 33 490
rect -33 416 33 432
rect -33 382 -17 416
rect 17 382 33 416
rect -33 366 33 382
rect -15 344 15 366
rect -15 238 15 260
rect -33 222 33 238
rect -33 188 -17 222
rect 17 188 33 222
rect -33 172 33 188
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -33 64 33 80
rect -15 42 15 64
rect -15 -64 15 -42
rect -33 -80 33 -64
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
rect -33 -188 33 -172
rect -33 -222 -17 -188
rect 17 -222 33 -188
rect -33 -238 33 -222
rect -15 -260 15 -238
rect -15 -366 15 -344
rect -33 -382 33 -366
rect -33 -416 -17 -382
rect 17 -416 33 -382
rect -33 -432 33 -416
rect -33 -490 33 -474
rect -33 -524 -17 -490
rect 17 -524 33 -490
rect -33 -540 33 -524
rect -15 -562 15 -540
rect -15 -668 15 -646
rect -33 -684 33 -668
rect -33 -718 -17 -684
rect 17 -718 33 -684
rect -33 -734 33 -718
rect -33 -792 33 -776
rect -33 -826 -17 -792
rect 17 -826 33 -792
rect -33 -842 33 -826
rect -15 -864 15 -842
rect -15 -970 15 -948
rect -33 -986 33 -970
rect -33 -1020 -17 -986
rect 17 -1020 33 -986
rect -33 -1036 33 -1020
<< polycont >>
rect -17 986 17 1020
rect -17 792 17 826
rect -17 684 17 718
rect -17 490 17 524
rect -17 382 17 416
rect -17 188 17 222
rect -17 80 17 114
rect -17 -114 17 -80
rect -17 -222 17 -188
rect -17 -416 17 -382
rect -17 -524 17 -490
rect -17 -718 17 -684
rect -17 -826 17 -792
rect -17 -1020 17 -986
<< locali >>
rect -175 1088 -79 1122
rect 79 1088 175 1122
rect -175 1026 -141 1088
rect 141 1026 175 1088
rect -33 986 -17 1020
rect 17 986 33 1020
rect -61 936 -27 952
rect -61 860 -27 876
rect 27 936 61 952
rect 27 860 61 876
rect -33 792 -17 826
rect 17 792 33 826
rect -33 684 -17 718
rect 17 684 33 718
rect -61 634 -27 650
rect -61 558 -27 574
rect 27 634 61 650
rect 27 558 61 574
rect -33 490 -17 524
rect 17 490 33 524
rect -33 382 -17 416
rect 17 382 33 416
rect -61 332 -27 348
rect -61 256 -27 272
rect 27 332 61 348
rect 27 256 61 272
rect -33 188 -17 222
rect 17 188 33 222
rect -33 80 -17 114
rect 17 80 33 114
rect -61 30 -27 46
rect -61 -46 -27 -30
rect 27 30 61 46
rect 27 -46 61 -30
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -222 -17 -188
rect 17 -222 33 -188
rect -61 -272 -27 -256
rect -61 -348 -27 -332
rect 27 -272 61 -256
rect 27 -348 61 -332
rect -33 -416 -17 -382
rect 17 -416 33 -382
rect -33 -524 -17 -490
rect 17 -524 33 -490
rect -61 -574 -27 -558
rect -61 -650 -27 -634
rect 27 -574 61 -558
rect 27 -650 61 -634
rect -33 -718 -17 -684
rect 17 -718 33 -684
rect -33 -826 -17 -792
rect 17 -826 33 -792
rect -61 -876 -27 -860
rect -61 -952 -27 -936
rect 27 -876 61 -860
rect 27 -952 61 -936
rect -33 -1020 -17 -986
rect 17 -1020 33 -986
rect -175 -1088 -141 -1026
rect 141 -1088 175 -1026
rect -175 -1122 -79 -1088
rect 79 -1122 175 -1088
<< viali >>
rect -17 986 17 1020
rect -61 876 -27 936
rect 27 876 61 936
rect -17 792 17 826
rect -17 684 17 718
rect -61 574 -27 634
rect 27 574 61 634
rect -17 490 17 524
rect -17 382 17 416
rect -61 272 -27 332
rect 27 272 61 332
rect -17 188 17 222
rect -17 80 17 114
rect -61 -30 -27 30
rect 27 -30 61 30
rect -17 -114 17 -80
rect -17 -222 17 -188
rect -61 -332 -27 -272
rect 27 -332 61 -272
rect -17 -416 17 -382
rect -17 -524 17 -490
rect -61 -634 -27 -574
rect 27 -634 61 -574
rect -17 -718 17 -684
rect -17 -826 17 -792
rect -61 -936 -27 -876
rect 27 -936 61 -876
rect -17 -1020 17 -986
<< metal1 >>
rect -29 1020 29 1026
rect -29 986 -17 1020
rect 17 986 29 1020
rect -29 980 29 986
rect -67 936 -21 948
rect -67 876 -61 936
rect -27 876 -21 936
rect -67 864 -21 876
rect 21 936 67 948
rect 21 876 27 936
rect 61 876 67 936
rect 21 864 67 876
rect -29 826 29 832
rect -29 792 -17 826
rect 17 792 29 826
rect -29 786 29 792
rect -29 718 29 724
rect -29 684 -17 718
rect 17 684 29 718
rect -29 678 29 684
rect -67 634 -21 646
rect -67 574 -61 634
rect -27 574 -21 634
rect -67 562 -21 574
rect 21 634 67 646
rect 21 574 27 634
rect 61 574 67 634
rect 21 562 67 574
rect -29 524 29 530
rect -29 490 -17 524
rect 17 490 29 524
rect -29 484 29 490
rect -29 416 29 422
rect -29 382 -17 416
rect 17 382 29 416
rect -29 376 29 382
rect -67 332 -21 344
rect -67 272 -61 332
rect -27 272 -21 332
rect -67 260 -21 272
rect 21 332 67 344
rect 21 272 27 332
rect 61 272 67 332
rect 21 260 67 272
rect -29 222 29 228
rect -29 188 -17 222
rect 17 188 29 222
rect -29 182 29 188
rect -29 114 29 120
rect -29 80 -17 114
rect 17 80 29 114
rect -29 74 29 80
rect -67 30 -21 42
rect -67 -30 -61 30
rect -27 -30 -21 30
rect -67 -42 -21 -30
rect 21 30 67 42
rect 21 -30 27 30
rect 61 -30 67 30
rect 21 -42 67 -30
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect -29 -120 29 -114
rect -29 -188 29 -182
rect -29 -222 -17 -188
rect 17 -222 29 -188
rect -29 -228 29 -222
rect -67 -272 -21 -260
rect -67 -332 -61 -272
rect -27 -332 -21 -272
rect -67 -344 -21 -332
rect 21 -272 67 -260
rect 21 -332 27 -272
rect 61 -332 67 -272
rect 21 -344 67 -332
rect -29 -382 29 -376
rect -29 -416 -17 -382
rect 17 -416 29 -382
rect -29 -422 29 -416
rect -29 -490 29 -484
rect -29 -524 -17 -490
rect 17 -524 29 -490
rect -29 -530 29 -524
rect -67 -574 -21 -562
rect -67 -634 -61 -574
rect -27 -634 -21 -574
rect -67 -646 -21 -634
rect 21 -574 67 -562
rect 21 -634 27 -574
rect 61 -634 67 -574
rect 21 -646 67 -634
rect -29 -684 29 -678
rect -29 -718 -17 -684
rect 17 -718 29 -684
rect -29 -724 29 -718
rect -29 -792 29 -786
rect -29 -826 -17 -792
rect 17 -826 29 -792
rect -29 -832 29 -826
rect -67 -876 -21 -864
rect -67 -936 -61 -876
rect -27 -936 -21 -876
rect -67 -948 -21 -936
rect 21 -876 67 -864
rect 21 -936 27 -876
rect 61 -936 67 -876
rect 21 -948 67 -936
rect -29 -986 29 -980
rect -29 -1020 -17 -986
rect 17 -1020 29 -986
rect -29 -1026 29 -1020
<< properties >>
string FIXED_BBOX -158 -1105 158 1105
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 7 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
