magic
tech sky130A
magscale 1 2
timestamp 1697806833
<< nwell >>
rect -28979 -3219 28979 3219
<< pmos >>
rect -28783 -3000 -26783 3000
rect -26725 -3000 -24725 3000
rect -24667 -3000 -22667 3000
rect -22609 -3000 -20609 3000
rect -20551 -3000 -18551 3000
rect -18493 -3000 -16493 3000
rect -16435 -3000 -14435 3000
rect -14377 -3000 -12377 3000
rect -12319 -3000 -10319 3000
rect -10261 -3000 -8261 3000
rect -8203 -3000 -6203 3000
rect -6145 -3000 -4145 3000
rect -4087 -3000 -2087 3000
rect -2029 -3000 -29 3000
rect 29 -3000 2029 3000
rect 2087 -3000 4087 3000
rect 4145 -3000 6145 3000
rect 6203 -3000 8203 3000
rect 8261 -3000 10261 3000
rect 10319 -3000 12319 3000
rect 12377 -3000 14377 3000
rect 14435 -3000 16435 3000
rect 16493 -3000 18493 3000
rect 18551 -3000 20551 3000
rect 20609 -3000 22609 3000
rect 22667 -3000 24667 3000
rect 24725 -3000 26725 3000
rect 26783 -3000 28783 3000
<< pdiff >>
rect -28841 2988 -28783 3000
rect -28841 -2988 -28829 2988
rect -28795 -2988 -28783 2988
rect -28841 -3000 -28783 -2988
rect -26783 2988 -26725 3000
rect -26783 -2988 -26771 2988
rect -26737 -2988 -26725 2988
rect -26783 -3000 -26725 -2988
rect -24725 2988 -24667 3000
rect -24725 -2988 -24713 2988
rect -24679 -2988 -24667 2988
rect -24725 -3000 -24667 -2988
rect -22667 2988 -22609 3000
rect -22667 -2988 -22655 2988
rect -22621 -2988 -22609 2988
rect -22667 -3000 -22609 -2988
rect -20609 2988 -20551 3000
rect -20609 -2988 -20597 2988
rect -20563 -2988 -20551 2988
rect -20609 -3000 -20551 -2988
rect -18551 2988 -18493 3000
rect -18551 -2988 -18539 2988
rect -18505 -2988 -18493 2988
rect -18551 -3000 -18493 -2988
rect -16493 2988 -16435 3000
rect -16493 -2988 -16481 2988
rect -16447 -2988 -16435 2988
rect -16493 -3000 -16435 -2988
rect -14435 2988 -14377 3000
rect -14435 -2988 -14423 2988
rect -14389 -2988 -14377 2988
rect -14435 -3000 -14377 -2988
rect -12377 2988 -12319 3000
rect -12377 -2988 -12365 2988
rect -12331 -2988 -12319 2988
rect -12377 -3000 -12319 -2988
rect -10319 2988 -10261 3000
rect -10319 -2988 -10307 2988
rect -10273 -2988 -10261 2988
rect -10319 -3000 -10261 -2988
rect -8261 2988 -8203 3000
rect -8261 -2988 -8249 2988
rect -8215 -2988 -8203 2988
rect -8261 -3000 -8203 -2988
rect -6203 2988 -6145 3000
rect -6203 -2988 -6191 2988
rect -6157 -2988 -6145 2988
rect -6203 -3000 -6145 -2988
rect -4145 2988 -4087 3000
rect -4145 -2988 -4133 2988
rect -4099 -2988 -4087 2988
rect -4145 -3000 -4087 -2988
rect -2087 2988 -2029 3000
rect -2087 -2988 -2075 2988
rect -2041 -2988 -2029 2988
rect -2087 -3000 -2029 -2988
rect -29 2988 29 3000
rect -29 -2988 -17 2988
rect 17 -2988 29 2988
rect -29 -3000 29 -2988
rect 2029 2988 2087 3000
rect 2029 -2988 2041 2988
rect 2075 -2988 2087 2988
rect 2029 -3000 2087 -2988
rect 4087 2988 4145 3000
rect 4087 -2988 4099 2988
rect 4133 -2988 4145 2988
rect 4087 -3000 4145 -2988
rect 6145 2988 6203 3000
rect 6145 -2988 6157 2988
rect 6191 -2988 6203 2988
rect 6145 -3000 6203 -2988
rect 8203 2988 8261 3000
rect 8203 -2988 8215 2988
rect 8249 -2988 8261 2988
rect 8203 -3000 8261 -2988
rect 10261 2988 10319 3000
rect 10261 -2988 10273 2988
rect 10307 -2988 10319 2988
rect 10261 -3000 10319 -2988
rect 12319 2988 12377 3000
rect 12319 -2988 12331 2988
rect 12365 -2988 12377 2988
rect 12319 -3000 12377 -2988
rect 14377 2988 14435 3000
rect 14377 -2988 14389 2988
rect 14423 -2988 14435 2988
rect 14377 -3000 14435 -2988
rect 16435 2988 16493 3000
rect 16435 -2988 16447 2988
rect 16481 -2988 16493 2988
rect 16435 -3000 16493 -2988
rect 18493 2988 18551 3000
rect 18493 -2988 18505 2988
rect 18539 -2988 18551 2988
rect 18493 -3000 18551 -2988
rect 20551 2988 20609 3000
rect 20551 -2988 20563 2988
rect 20597 -2988 20609 2988
rect 20551 -3000 20609 -2988
rect 22609 2988 22667 3000
rect 22609 -2988 22621 2988
rect 22655 -2988 22667 2988
rect 22609 -3000 22667 -2988
rect 24667 2988 24725 3000
rect 24667 -2988 24679 2988
rect 24713 -2988 24725 2988
rect 24667 -3000 24725 -2988
rect 26725 2988 26783 3000
rect 26725 -2988 26737 2988
rect 26771 -2988 26783 2988
rect 26725 -3000 26783 -2988
rect 28783 2988 28841 3000
rect 28783 -2988 28795 2988
rect 28829 -2988 28841 2988
rect 28783 -3000 28841 -2988
<< pdiffc >>
rect -28829 -2988 -28795 2988
rect -26771 -2988 -26737 2988
rect -24713 -2988 -24679 2988
rect -22655 -2988 -22621 2988
rect -20597 -2988 -20563 2988
rect -18539 -2988 -18505 2988
rect -16481 -2988 -16447 2988
rect -14423 -2988 -14389 2988
rect -12365 -2988 -12331 2988
rect -10307 -2988 -10273 2988
rect -8249 -2988 -8215 2988
rect -6191 -2988 -6157 2988
rect -4133 -2988 -4099 2988
rect -2075 -2988 -2041 2988
rect -17 -2988 17 2988
rect 2041 -2988 2075 2988
rect 4099 -2988 4133 2988
rect 6157 -2988 6191 2988
rect 8215 -2988 8249 2988
rect 10273 -2988 10307 2988
rect 12331 -2988 12365 2988
rect 14389 -2988 14423 2988
rect 16447 -2988 16481 2988
rect 18505 -2988 18539 2988
rect 20563 -2988 20597 2988
rect 22621 -2988 22655 2988
rect 24679 -2988 24713 2988
rect 26737 -2988 26771 2988
rect 28795 -2988 28829 2988
<< nsubdiff >>
rect -28943 3149 -28847 3183
rect 28847 3149 28943 3183
rect -28943 3087 -28909 3149
rect 28909 3087 28943 3149
rect -28943 -3149 -28909 -3087
rect 28909 -3149 28943 -3087
rect -28943 -3183 -28847 -3149
rect 28847 -3183 28943 -3149
<< nsubdiffcont >>
rect -28847 3149 28847 3183
rect -28943 -3087 -28909 3087
rect 28909 -3087 28943 3087
rect -28847 -3183 28847 -3149
<< poly >>
rect -28783 3081 -26783 3097
rect -28783 3047 -28767 3081
rect -26799 3047 -26783 3081
rect -28783 3000 -26783 3047
rect -26725 3081 -24725 3097
rect -26725 3047 -26709 3081
rect -24741 3047 -24725 3081
rect -26725 3000 -24725 3047
rect -24667 3081 -22667 3097
rect -24667 3047 -24651 3081
rect -22683 3047 -22667 3081
rect -24667 3000 -22667 3047
rect -22609 3081 -20609 3097
rect -22609 3047 -22593 3081
rect -20625 3047 -20609 3081
rect -22609 3000 -20609 3047
rect -20551 3081 -18551 3097
rect -20551 3047 -20535 3081
rect -18567 3047 -18551 3081
rect -20551 3000 -18551 3047
rect -18493 3081 -16493 3097
rect -18493 3047 -18477 3081
rect -16509 3047 -16493 3081
rect -18493 3000 -16493 3047
rect -16435 3081 -14435 3097
rect -16435 3047 -16419 3081
rect -14451 3047 -14435 3081
rect -16435 3000 -14435 3047
rect -14377 3081 -12377 3097
rect -14377 3047 -14361 3081
rect -12393 3047 -12377 3081
rect -14377 3000 -12377 3047
rect -12319 3081 -10319 3097
rect -12319 3047 -12303 3081
rect -10335 3047 -10319 3081
rect -12319 3000 -10319 3047
rect -10261 3081 -8261 3097
rect -10261 3047 -10245 3081
rect -8277 3047 -8261 3081
rect -10261 3000 -8261 3047
rect -8203 3081 -6203 3097
rect -8203 3047 -8187 3081
rect -6219 3047 -6203 3081
rect -8203 3000 -6203 3047
rect -6145 3081 -4145 3097
rect -6145 3047 -6129 3081
rect -4161 3047 -4145 3081
rect -6145 3000 -4145 3047
rect -4087 3081 -2087 3097
rect -4087 3047 -4071 3081
rect -2103 3047 -2087 3081
rect -4087 3000 -2087 3047
rect -2029 3081 -29 3097
rect -2029 3047 -2013 3081
rect -45 3047 -29 3081
rect -2029 3000 -29 3047
rect 29 3081 2029 3097
rect 29 3047 45 3081
rect 2013 3047 2029 3081
rect 29 3000 2029 3047
rect 2087 3081 4087 3097
rect 2087 3047 2103 3081
rect 4071 3047 4087 3081
rect 2087 3000 4087 3047
rect 4145 3081 6145 3097
rect 4145 3047 4161 3081
rect 6129 3047 6145 3081
rect 4145 3000 6145 3047
rect 6203 3081 8203 3097
rect 6203 3047 6219 3081
rect 8187 3047 8203 3081
rect 6203 3000 8203 3047
rect 8261 3081 10261 3097
rect 8261 3047 8277 3081
rect 10245 3047 10261 3081
rect 8261 3000 10261 3047
rect 10319 3081 12319 3097
rect 10319 3047 10335 3081
rect 12303 3047 12319 3081
rect 10319 3000 12319 3047
rect 12377 3081 14377 3097
rect 12377 3047 12393 3081
rect 14361 3047 14377 3081
rect 12377 3000 14377 3047
rect 14435 3081 16435 3097
rect 14435 3047 14451 3081
rect 16419 3047 16435 3081
rect 14435 3000 16435 3047
rect 16493 3081 18493 3097
rect 16493 3047 16509 3081
rect 18477 3047 18493 3081
rect 16493 3000 18493 3047
rect 18551 3081 20551 3097
rect 18551 3047 18567 3081
rect 20535 3047 20551 3081
rect 18551 3000 20551 3047
rect 20609 3081 22609 3097
rect 20609 3047 20625 3081
rect 22593 3047 22609 3081
rect 20609 3000 22609 3047
rect 22667 3081 24667 3097
rect 22667 3047 22683 3081
rect 24651 3047 24667 3081
rect 22667 3000 24667 3047
rect 24725 3081 26725 3097
rect 24725 3047 24741 3081
rect 26709 3047 26725 3081
rect 24725 3000 26725 3047
rect 26783 3081 28783 3097
rect 26783 3047 26799 3081
rect 28767 3047 28783 3081
rect 26783 3000 28783 3047
rect -28783 -3047 -26783 -3000
rect -28783 -3081 -28767 -3047
rect -26799 -3081 -26783 -3047
rect -28783 -3097 -26783 -3081
rect -26725 -3047 -24725 -3000
rect -26725 -3081 -26709 -3047
rect -24741 -3081 -24725 -3047
rect -26725 -3097 -24725 -3081
rect -24667 -3047 -22667 -3000
rect -24667 -3081 -24651 -3047
rect -22683 -3081 -22667 -3047
rect -24667 -3097 -22667 -3081
rect -22609 -3047 -20609 -3000
rect -22609 -3081 -22593 -3047
rect -20625 -3081 -20609 -3047
rect -22609 -3097 -20609 -3081
rect -20551 -3047 -18551 -3000
rect -20551 -3081 -20535 -3047
rect -18567 -3081 -18551 -3047
rect -20551 -3097 -18551 -3081
rect -18493 -3047 -16493 -3000
rect -18493 -3081 -18477 -3047
rect -16509 -3081 -16493 -3047
rect -18493 -3097 -16493 -3081
rect -16435 -3047 -14435 -3000
rect -16435 -3081 -16419 -3047
rect -14451 -3081 -14435 -3047
rect -16435 -3097 -14435 -3081
rect -14377 -3047 -12377 -3000
rect -14377 -3081 -14361 -3047
rect -12393 -3081 -12377 -3047
rect -14377 -3097 -12377 -3081
rect -12319 -3047 -10319 -3000
rect -12319 -3081 -12303 -3047
rect -10335 -3081 -10319 -3047
rect -12319 -3097 -10319 -3081
rect -10261 -3047 -8261 -3000
rect -10261 -3081 -10245 -3047
rect -8277 -3081 -8261 -3047
rect -10261 -3097 -8261 -3081
rect -8203 -3047 -6203 -3000
rect -8203 -3081 -8187 -3047
rect -6219 -3081 -6203 -3047
rect -8203 -3097 -6203 -3081
rect -6145 -3047 -4145 -3000
rect -6145 -3081 -6129 -3047
rect -4161 -3081 -4145 -3047
rect -6145 -3097 -4145 -3081
rect -4087 -3047 -2087 -3000
rect -4087 -3081 -4071 -3047
rect -2103 -3081 -2087 -3047
rect -4087 -3097 -2087 -3081
rect -2029 -3047 -29 -3000
rect -2029 -3081 -2013 -3047
rect -45 -3081 -29 -3047
rect -2029 -3097 -29 -3081
rect 29 -3047 2029 -3000
rect 29 -3081 45 -3047
rect 2013 -3081 2029 -3047
rect 29 -3097 2029 -3081
rect 2087 -3047 4087 -3000
rect 2087 -3081 2103 -3047
rect 4071 -3081 4087 -3047
rect 2087 -3097 4087 -3081
rect 4145 -3047 6145 -3000
rect 4145 -3081 4161 -3047
rect 6129 -3081 6145 -3047
rect 4145 -3097 6145 -3081
rect 6203 -3047 8203 -3000
rect 6203 -3081 6219 -3047
rect 8187 -3081 8203 -3047
rect 6203 -3097 8203 -3081
rect 8261 -3047 10261 -3000
rect 8261 -3081 8277 -3047
rect 10245 -3081 10261 -3047
rect 8261 -3097 10261 -3081
rect 10319 -3047 12319 -3000
rect 10319 -3081 10335 -3047
rect 12303 -3081 12319 -3047
rect 10319 -3097 12319 -3081
rect 12377 -3047 14377 -3000
rect 12377 -3081 12393 -3047
rect 14361 -3081 14377 -3047
rect 12377 -3097 14377 -3081
rect 14435 -3047 16435 -3000
rect 14435 -3081 14451 -3047
rect 16419 -3081 16435 -3047
rect 14435 -3097 16435 -3081
rect 16493 -3047 18493 -3000
rect 16493 -3081 16509 -3047
rect 18477 -3081 18493 -3047
rect 16493 -3097 18493 -3081
rect 18551 -3047 20551 -3000
rect 18551 -3081 18567 -3047
rect 20535 -3081 20551 -3047
rect 18551 -3097 20551 -3081
rect 20609 -3047 22609 -3000
rect 20609 -3081 20625 -3047
rect 22593 -3081 22609 -3047
rect 20609 -3097 22609 -3081
rect 22667 -3047 24667 -3000
rect 22667 -3081 22683 -3047
rect 24651 -3081 24667 -3047
rect 22667 -3097 24667 -3081
rect 24725 -3047 26725 -3000
rect 24725 -3081 24741 -3047
rect 26709 -3081 26725 -3047
rect 24725 -3097 26725 -3081
rect 26783 -3047 28783 -3000
rect 26783 -3081 26799 -3047
rect 28767 -3081 28783 -3047
rect 26783 -3097 28783 -3081
<< polycont >>
rect -28767 3047 -26799 3081
rect -26709 3047 -24741 3081
rect -24651 3047 -22683 3081
rect -22593 3047 -20625 3081
rect -20535 3047 -18567 3081
rect -18477 3047 -16509 3081
rect -16419 3047 -14451 3081
rect -14361 3047 -12393 3081
rect -12303 3047 -10335 3081
rect -10245 3047 -8277 3081
rect -8187 3047 -6219 3081
rect -6129 3047 -4161 3081
rect -4071 3047 -2103 3081
rect -2013 3047 -45 3081
rect 45 3047 2013 3081
rect 2103 3047 4071 3081
rect 4161 3047 6129 3081
rect 6219 3047 8187 3081
rect 8277 3047 10245 3081
rect 10335 3047 12303 3081
rect 12393 3047 14361 3081
rect 14451 3047 16419 3081
rect 16509 3047 18477 3081
rect 18567 3047 20535 3081
rect 20625 3047 22593 3081
rect 22683 3047 24651 3081
rect 24741 3047 26709 3081
rect 26799 3047 28767 3081
rect -28767 -3081 -26799 -3047
rect -26709 -3081 -24741 -3047
rect -24651 -3081 -22683 -3047
rect -22593 -3081 -20625 -3047
rect -20535 -3081 -18567 -3047
rect -18477 -3081 -16509 -3047
rect -16419 -3081 -14451 -3047
rect -14361 -3081 -12393 -3047
rect -12303 -3081 -10335 -3047
rect -10245 -3081 -8277 -3047
rect -8187 -3081 -6219 -3047
rect -6129 -3081 -4161 -3047
rect -4071 -3081 -2103 -3047
rect -2013 -3081 -45 -3047
rect 45 -3081 2013 -3047
rect 2103 -3081 4071 -3047
rect 4161 -3081 6129 -3047
rect 6219 -3081 8187 -3047
rect 8277 -3081 10245 -3047
rect 10335 -3081 12303 -3047
rect 12393 -3081 14361 -3047
rect 14451 -3081 16419 -3047
rect 16509 -3081 18477 -3047
rect 18567 -3081 20535 -3047
rect 20625 -3081 22593 -3047
rect 22683 -3081 24651 -3047
rect 24741 -3081 26709 -3047
rect 26799 -3081 28767 -3047
<< locali >>
rect -28943 3149 -28847 3183
rect 28847 3149 28943 3183
rect -28943 3087 -28909 3149
rect 28909 3087 28943 3149
rect -28783 3047 -28767 3081
rect -26799 3047 -26783 3081
rect -26725 3047 -26709 3081
rect -24741 3047 -24725 3081
rect -24667 3047 -24651 3081
rect -22683 3047 -22667 3081
rect -22609 3047 -22593 3081
rect -20625 3047 -20609 3081
rect -20551 3047 -20535 3081
rect -18567 3047 -18551 3081
rect -18493 3047 -18477 3081
rect -16509 3047 -16493 3081
rect -16435 3047 -16419 3081
rect -14451 3047 -14435 3081
rect -14377 3047 -14361 3081
rect -12393 3047 -12377 3081
rect -12319 3047 -12303 3081
rect -10335 3047 -10319 3081
rect -10261 3047 -10245 3081
rect -8277 3047 -8261 3081
rect -8203 3047 -8187 3081
rect -6219 3047 -6203 3081
rect -6145 3047 -6129 3081
rect -4161 3047 -4145 3081
rect -4087 3047 -4071 3081
rect -2103 3047 -2087 3081
rect -2029 3047 -2013 3081
rect -45 3047 -29 3081
rect 29 3047 45 3081
rect 2013 3047 2029 3081
rect 2087 3047 2103 3081
rect 4071 3047 4087 3081
rect 4145 3047 4161 3081
rect 6129 3047 6145 3081
rect 6203 3047 6219 3081
rect 8187 3047 8203 3081
rect 8261 3047 8277 3081
rect 10245 3047 10261 3081
rect 10319 3047 10335 3081
rect 12303 3047 12319 3081
rect 12377 3047 12393 3081
rect 14361 3047 14377 3081
rect 14435 3047 14451 3081
rect 16419 3047 16435 3081
rect 16493 3047 16509 3081
rect 18477 3047 18493 3081
rect 18551 3047 18567 3081
rect 20535 3047 20551 3081
rect 20609 3047 20625 3081
rect 22593 3047 22609 3081
rect 22667 3047 22683 3081
rect 24651 3047 24667 3081
rect 24725 3047 24741 3081
rect 26709 3047 26725 3081
rect 26783 3047 26799 3081
rect 28767 3047 28783 3081
rect -28829 2988 -28795 3004
rect -28829 -3004 -28795 -2988
rect -26771 2988 -26737 3004
rect -26771 -3004 -26737 -2988
rect -24713 2988 -24679 3004
rect -24713 -3004 -24679 -2988
rect -22655 2988 -22621 3004
rect -22655 -3004 -22621 -2988
rect -20597 2988 -20563 3004
rect -20597 -3004 -20563 -2988
rect -18539 2988 -18505 3004
rect -18539 -3004 -18505 -2988
rect -16481 2988 -16447 3004
rect -16481 -3004 -16447 -2988
rect -14423 2988 -14389 3004
rect -14423 -3004 -14389 -2988
rect -12365 2988 -12331 3004
rect -12365 -3004 -12331 -2988
rect -10307 2988 -10273 3004
rect -10307 -3004 -10273 -2988
rect -8249 2988 -8215 3004
rect -8249 -3004 -8215 -2988
rect -6191 2988 -6157 3004
rect -6191 -3004 -6157 -2988
rect -4133 2988 -4099 3004
rect -4133 -3004 -4099 -2988
rect -2075 2988 -2041 3004
rect -2075 -3004 -2041 -2988
rect -17 2988 17 3004
rect -17 -3004 17 -2988
rect 2041 2988 2075 3004
rect 2041 -3004 2075 -2988
rect 4099 2988 4133 3004
rect 4099 -3004 4133 -2988
rect 6157 2988 6191 3004
rect 6157 -3004 6191 -2988
rect 8215 2988 8249 3004
rect 8215 -3004 8249 -2988
rect 10273 2988 10307 3004
rect 10273 -3004 10307 -2988
rect 12331 2988 12365 3004
rect 12331 -3004 12365 -2988
rect 14389 2988 14423 3004
rect 14389 -3004 14423 -2988
rect 16447 2988 16481 3004
rect 16447 -3004 16481 -2988
rect 18505 2988 18539 3004
rect 18505 -3004 18539 -2988
rect 20563 2988 20597 3004
rect 20563 -3004 20597 -2988
rect 22621 2988 22655 3004
rect 22621 -3004 22655 -2988
rect 24679 2988 24713 3004
rect 24679 -3004 24713 -2988
rect 26737 2988 26771 3004
rect 26737 -3004 26771 -2988
rect 28795 2988 28829 3004
rect 28795 -3004 28829 -2988
rect -28783 -3081 -28767 -3047
rect -26799 -3081 -26783 -3047
rect -26725 -3081 -26709 -3047
rect -24741 -3081 -24725 -3047
rect -24667 -3081 -24651 -3047
rect -22683 -3081 -22667 -3047
rect -22609 -3081 -22593 -3047
rect -20625 -3081 -20609 -3047
rect -20551 -3081 -20535 -3047
rect -18567 -3081 -18551 -3047
rect -18493 -3081 -18477 -3047
rect -16509 -3081 -16493 -3047
rect -16435 -3081 -16419 -3047
rect -14451 -3081 -14435 -3047
rect -14377 -3081 -14361 -3047
rect -12393 -3081 -12377 -3047
rect -12319 -3081 -12303 -3047
rect -10335 -3081 -10319 -3047
rect -10261 -3081 -10245 -3047
rect -8277 -3081 -8261 -3047
rect -8203 -3081 -8187 -3047
rect -6219 -3081 -6203 -3047
rect -6145 -3081 -6129 -3047
rect -4161 -3081 -4145 -3047
rect -4087 -3081 -4071 -3047
rect -2103 -3081 -2087 -3047
rect -2029 -3081 -2013 -3047
rect -45 -3081 -29 -3047
rect 29 -3081 45 -3047
rect 2013 -3081 2029 -3047
rect 2087 -3081 2103 -3047
rect 4071 -3081 4087 -3047
rect 4145 -3081 4161 -3047
rect 6129 -3081 6145 -3047
rect 6203 -3081 6219 -3047
rect 8187 -3081 8203 -3047
rect 8261 -3081 8277 -3047
rect 10245 -3081 10261 -3047
rect 10319 -3081 10335 -3047
rect 12303 -3081 12319 -3047
rect 12377 -3081 12393 -3047
rect 14361 -3081 14377 -3047
rect 14435 -3081 14451 -3047
rect 16419 -3081 16435 -3047
rect 16493 -3081 16509 -3047
rect 18477 -3081 18493 -3047
rect 18551 -3081 18567 -3047
rect 20535 -3081 20551 -3047
rect 20609 -3081 20625 -3047
rect 22593 -3081 22609 -3047
rect 22667 -3081 22683 -3047
rect 24651 -3081 24667 -3047
rect 24725 -3081 24741 -3047
rect 26709 -3081 26725 -3047
rect 26783 -3081 26799 -3047
rect 28767 -3081 28783 -3047
rect -28943 -3149 -28909 -3087
rect 28909 -3149 28943 -3087
rect -28943 -3183 -28847 -3149
rect 28847 -3183 28943 -3149
<< viali >>
rect -28767 3047 -26799 3081
rect -26709 3047 -24741 3081
rect -24651 3047 -22683 3081
rect -22593 3047 -20625 3081
rect -20535 3047 -18567 3081
rect -18477 3047 -16509 3081
rect -16419 3047 -14451 3081
rect -14361 3047 -12393 3081
rect -12303 3047 -10335 3081
rect -10245 3047 -8277 3081
rect -8187 3047 -6219 3081
rect -6129 3047 -4161 3081
rect -4071 3047 -2103 3081
rect -2013 3047 -45 3081
rect 45 3047 2013 3081
rect 2103 3047 4071 3081
rect 4161 3047 6129 3081
rect 6219 3047 8187 3081
rect 8277 3047 10245 3081
rect 10335 3047 12303 3081
rect 12393 3047 14361 3081
rect 14451 3047 16419 3081
rect 16509 3047 18477 3081
rect 18567 3047 20535 3081
rect 20625 3047 22593 3081
rect 22683 3047 24651 3081
rect 24741 3047 26709 3081
rect 26799 3047 28767 3081
rect -28829 -2988 -28795 2988
rect -26771 -2988 -26737 2988
rect -24713 -2988 -24679 2988
rect -22655 -2988 -22621 2988
rect -20597 -2988 -20563 2988
rect -18539 -2988 -18505 2988
rect -16481 -2988 -16447 2988
rect -14423 -2988 -14389 2988
rect -12365 -2988 -12331 2988
rect -10307 -2988 -10273 2988
rect -8249 -2988 -8215 2988
rect -6191 -2988 -6157 2988
rect -4133 -2988 -4099 2988
rect -2075 -2988 -2041 2988
rect -17 -2988 17 2988
rect 2041 -2988 2075 2988
rect 4099 -2988 4133 2988
rect 6157 -2988 6191 2988
rect 8215 -2988 8249 2988
rect 10273 -2988 10307 2988
rect 12331 -2988 12365 2988
rect 14389 -2988 14423 2988
rect 16447 -2988 16481 2988
rect 18505 -2988 18539 2988
rect 20563 -2988 20597 2988
rect 22621 -2988 22655 2988
rect 24679 -2988 24713 2988
rect 26737 -2988 26771 2988
rect 28795 -2988 28829 2988
rect -28767 -3081 -26799 -3047
rect -26709 -3081 -24741 -3047
rect -24651 -3081 -22683 -3047
rect -22593 -3081 -20625 -3047
rect -20535 -3081 -18567 -3047
rect -18477 -3081 -16509 -3047
rect -16419 -3081 -14451 -3047
rect -14361 -3081 -12393 -3047
rect -12303 -3081 -10335 -3047
rect -10245 -3081 -8277 -3047
rect -8187 -3081 -6219 -3047
rect -6129 -3081 -4161 -3047
rect -4071 -3081 -2103 -3047
rect -2013 -3081 -45 -3047
rect 45 -3081 2013 -3047
rect 2103 -3081 4071 -3047
rect 4161 -3081 6129 -3047
rect 6219 -3081 8187 -3047
rect 8277 -3081 10245 -3047
rect 10335 -3081 12303 -3047
rect 12393 -3081 14361 -3047
rect 14451 -3081 16419 -3047
rect 16509 -3081 18477 -3047
rect 18567 -3081 20535 -3047
rect 20625 -3081 22593 -3047
rect 22683 -3081 24651 -3047
rect 24741 -3081 26709 -3047
rect 26799 -3081 28767 -3047
<< metal1 >>
rect -28779 3081 -26787 3087
rect -28779 3047 -28767 3081
rect -26799 3047 -26787 3081
rect -28779 3041 -26787 3047
rect -26721 3081 -24729 3087
rect -26721 3047 -26709 3081
rect -24741 3047 -24729 3081
rect -26721 3041 -24729 3047
rect -24663 3081 -22671 3087
rect -24663 3047 -24651 3081
rect -22683 3047 -22671 3081
rect -24663 3041 -22671 3047
rect -22605 3081 -20613 3087
rect -22605 3047 -22593 3081
rect -20625 3047 -20613 3081
rect -22605 3041 -20613 3047
rect -20547 3081 -18555 3087
rect -20547 3047 -20535 3081
rect -18567 3047 -18555 3081
rect -20547 3041 -18555 3047
rect -18489 3081 -16497 3087
rect -18489 3047 -18477 3081
rect -16509 3047 -16497 3081
rect -18489 3041 -16497 3047
rect -16431 3081 -14439 3087
rect -16431 3047 -16419 3081
rect -14451 3047 -14439 3081
rect -16431 3041 -14439 3047
rect -14373 3081 -12381 3087
rect -14373 3047 -14361 3081
rect -12393 3047 -12381 3081
rect -14373 3041 -12381 3047
rect -12315 3081 -10323 3087
rect -12315 3047 -12303 3081
rect -10335 3047 -10323 3081
rect -12315 3041 -10323 3047
rect -10257 3081 -8265 3087
rect -10257 3047 -10245 3081
rect -8277 3047 -8265 3081
rect -10257 3041 -8265 3047
rect -8199 3081 -6207 3087
rect -8199 3047 -8187 3081
rect -6219 3047 -6207 3081
rect -8199 3041 -6207 3047
rect -6141 3081 -4149 3087
rect -6141 3047 -6129 3081
rect -4161 3047 -4149 3081
rect -6141 3041 -4149 3047
rect -4083 3081 -2091 3087
rect -4083 3047 -4071 3081
rect -2103 3047 -2091 3081
rect -4083 3041 -2091 3047
rect -2025 3081 -33 3087
rect -2025 3047 -2013 3081
rect -45 3047 -33 3081
rect -2025 3041 -33 3047
rect 33 3081 2025 3087
rect 33 3047 45 3081
rect 2013 3047 2025 3081
rect 33 3041 2025 3047
rect 2091 3081 4083 3087
rect 2091 3047 2103 3081
rect 4071 3047 4083 3081
rect 2091 3041 4083 3047
rect 4149 3081 6141 3087
rect 4149 3047 4161 3081
rect 6129 3047 6141 3081
rect 4149 3041 6141 3047
rect 6207 3081 8199 3087
rect 6207 3047 6219 3081
rect 8187 3047 8199 3081
rect 6207 3041 8199 3047
rect 8265 3081 10257 3087
rect 8265 3047 8277 3081
rect 10245 3047 10257 3081
rect 8265 3041 10257 3047
rect 10323 3081 12315 3087
rect 10323 3047 10335 3081
rect 12303 3047 12315 3081
rect 10323 3041 12315 3047
rect 12381 3081 14373 3087
rect 12381 3047 12393 3081
rect 14361 3047 14373 3081
rect 12381 3041 14373 3047
rect 14439 3081 16431 3087
rect 14439 3047 14451 3081
rect 16419 3047 16431 3081
rect 14439 3041 16431 3047
rect 16497 3081 18489 3087
rect 16497 3047 16509 3081
rect 18477 3047 18489 3081
rect 16497 3041 18489 3047
rect 18555 3081 20547 3087
rect 18555 3047 18567 3081
rect 20535 3047 20547 3081
rect 18555 3041 20547 3047
rect 20613 3081 22605 3087
rect 20613 3047 20625 3081
rect 22593 3047 22605 3081
rect 20613 3041 22605 3047
rect 22671 3081 24663 3087
rect 22671 3047 22683 3081
rect 24651 3047 24663 3081
rect 22671 3041 24663 3047
rect 24729 3081 26721 3087
rect 24729 3047 24741 3081
rect 26709 3047 26721 3081
rect 24729 3041 26721 3047
rect 26787 3081 28779 3087
rect 26787 3047 26799 3081
rect 28767 3047 28779 3081
rect 26787 3041 28779 3047
rect -28835 2988 -28789 3000
rect -28835 -2988 -28829 2988
rect -28795 -2988 -28789 2988
rect -28835 -3000 -28789 -2988
rect -26777 2988 -26731 3000
rect -26777 -2988 -26771 2988
rect -26737 -2988 -26731 2988
rect -26777 -3000 -26731 -2988
rect -24719 2988 -24673 3000
rect -24719 -2988 -24713 2988
rect -24679 -2988 -24673 2988
rect -24719 -3000 -24673 -2988
rect -22661 2988 -22615 3000
rect -22661 -2988 -22655 2988
rect -22621 -2988 -22615 2988
rect -22661 -3000 -22615 -2988
rect -20603 2988 -20557 3000
rect -20603 -2988 -20597 2988
rect -20563 -2988 -20557 2988
rect -20603 -3000 -20557 -2988
rect -18545 2988 -18499 3000
rect -18545 -2988 -18539 2988
rect -18505 -2988 -18499 2988
rect -18545 -3000 -18499 -2988
rect -16487 2988 -16441 3000
rect -16487 -2988 -16481 2988
rect -16447 -2988 -16441 2988
rect -16487 -3000 -16441 -2988
rect -14429 2988 -14383 3000
rect -14429 -2988 -14423 2988
rect -14389 -2988 -14383 2988
rect -14429 -3000 -14383 -2988
rect -12371 2988 -12325 3000
rect -12371 -2988 -12365 2988
rect -12331 -2988 -12325 2988
rect -12371 -3000 -12325 -2988
rect -10313 2988 -10267 3000
rect -10313 -2988 -10307 2988
rect -10273 -2988 -10267 2988
rect -10313 -3000 -10267 -2988
rect -8255 2988 -8209 3000
rect -8255 -2988 -8249 2988
rect -8215 -2988 -8209 2988
rect -8255 -3000 -8209 -2988
rect -6197 2988 -6151 3000
rect -6197 -2988 -6191 2988
rect -6157 -2988 -6151 2988
rect -6197 -3000 -6151 -2988
rect -4139 2988 -4093 3000
rect -4139 -2988 -4133 2988
rect -4099 -2988 -4093 2988
rect -4139 -3000 -4093 -2988
rect -2081 2988 -2035 3000
rect -2081 -2988 -2075 2988
rect -2041 -2988 -2035 2988
rect -2081 -3000 -2035 -2988
rect -23 2988 23 3000
rect -23 -2988 -17 2988
rect 17 -2988 23 2988
rect -23 -3000 23 -2988
rect 2035 2988 2081 3000
rect 2035 -2988 2041 2988
rect 2075 -2988 2081 2988
rect 2035 -3000 2081 -2988
rect 4093 2988 4139 3000
rect 4093 -2988 4099 2988
rect 4133 -2988 4139 2988
rect 4093 -3000 4139 -2988
rect 6151 2988 6197 3000
rect 6151 -2988 6157 2988
rect 6191 -2988 6197 2988
rect 6151 -3000 6197 -2988
rect 8209 2988 8255 3000
rect 8209 -2988 8215 2988
rect 8249 -2988 8255 2988
rect 8209 -3000 8255 -2988
rect 10267 2988 10313 3000
rect 10267 -2988 10273 2988
rect 10307 -2988 10313 2988
rect 10267 -3000 10313 -2988
rect 12325 2988 12371 3000
rect 12325 -2988 12331 2988
rect 12365 -2988 12371 2988
rect 12325 -3000 12371 -2988
rect 14383 2988 14429 3000
rect 14383 -2988 14389 2988
rect 14423 -2988 14429 2988
rect 14383 -3000 14429 -2988
rect 16441 2988 16487 3000
rect 16441 -2988 16447 2988
rect 16481 -2988 16487 2988
rect 16441 -3000 16487 -2988
rect 18499 2988 18545 3000
rect 18499 -2988 18505 2988
rect 18539 -2988 18545 2988
rect 18499 -3000 18545 -2988
rect 20557 2988 20603 3000
rect 20557 -2988 20563 2988
rect 20597 -2988 20603 2988
rect 20557 -3000 20603 -2988
rect 22615 2988 22661 3000
rect 22615 -2988 22621 2988
rect 22655 -2988 22661 2988
rect 22615 -3000 22661 -2988
rect 24673 2988 24719 3000
rect 24673 -2988 24679 2988
rect 24713 -2988 24719 2988
rect 24673 -3000 24719 -2988
rect 26731 2988 26777 3000
rect 26731 -2988 26737 2988
rect 26771 -2988 26777 2988
rect 26731 -3000 26777 -2988
rect 28789 2988 28835 3000
rect 28789 -2988 28795 2988
rect 28829 -2988 28835 2988
rect 28789 -3000 28835 -2988
rect -28779 -3047 -26787 -3041
rect -28779 -3081 -28767 -3047
rect -26799 -3081 -26787 -3047
rect -28779 -3087 -26787 -3081
rect -26721 -3047 -24729 -3041
rect -26721 -3081 -26709 -3047
rect -24741 -3081 -24729 -3047
rect -26721 -3087 -24729 -3081
rect -24663 -3047 -22671 -3041
rect -24663 -3081 -24651 -3047
rect -22683 -3081 -22671 -3047
rect -24663 -3087 -22671 -3081
rect -22605 -3047 -20613 -3041
rect -22605 -3081 -22593 -3047
rect -20625 -3081 -20613 -3047
rect -22605 -3087 -20613 -3081
rect -20547 -3047 -18555 -3041
rect -20547 -3081 -20535 -3047
rect -18567 -3081 -18555 -3047
rect -20547 -3087 -18555 -3081
rect -18489 -3047 -16497 -3041
rect -18489 -3081 -18477 -3047
rect -16509 -3081 -16497 -3047
rect -18489 -3087 -16497 -3081
rect -16431 -3047 -14439 -3041
rect -16431 -3081 -16419 -3047
rect -14451 -3081 -14439 -3047
rect -16431 -3087 -14439 -3081
rect -14373 -3047 -12381 -3041
rect -14373 -3081 -14361 -3047
rect -12393 -3081 -12381 -3047
rect -14373 -3087 -12381 -3081
rect -12315 -3047 -10323 -3041
rect -12315 -3081 -12303 -3047
rect -10335 -3081 -10323 -3047
rect -12315 -3087 -10323 -3081
rect -10257 -3047 -8265 -3041
rect -10257 -3081 -10245 -3047
rect -8277 -3081 -8265 -3047
rect -10257 -3087 -8265 -3081
rect -8199 -3047 -6207 -3041
rect -8199 -3081 -8187 -3047
rect -6219 -3081 -6207 -3047
rect -8199 -3087 -6207 -3081
rect -6141 -3047 -4149 -3041
rect -6141 -3081 -6129 -3047
rect -4161 -3081 -4149 -3047
rect -6141 -3087 -4149 -3081
rect -4083 -3047 -2091 -3041
rect -4083 -3081 -4071 -3047
rect -2103 -3081 -2091 -3047
rect -4083 -3087 -2091 -3081
rect -2025 -3047 -33 -3041
rect -2025 -3081 -2013 -3047
rect -45 -3081 -33 -3047
rect -2025 -3087 -33 -3081
rect 33 -3047 2025 -3041
rect 33 -3081 45 -3047
rect 2013 -3081 2025 -3047
rect 33 -3087 2025 -3081
rect 2091 -3047 4083 -3041
rect 2091 -3081 2103 -3047
rect 4071 -3081 4083 -3047
rect 2091 -3087 4083 -3081
rect 4149 -3047 6141 -3041
rect 4149 -3081 4161 -3047
rect 6129 -3081 6141 -3047
rect 4149 -3087 6141 -3081
rect 6207 -3047 8199 -3041
rect 6207 -3081 6219 -3047
rect 8187 -3081 8199 -3047
rect 6207 -3087 8199 -3081
rect 8265 -3047 10257 -3041
rect 8265 -3081 8277 -3047
rect 10245 -3081 10257 -3047
rect 8265 -3087 10257 -3081
rect 10323 -3047 12315 -3041
rect 10323 -3081 10335 -3047
rect 12303 -3081 12315 -3047
rect 10323 -3087 12315 -3081
rect 12381 -3047 14373 -3041
rect 12381 -3081 12393 -3047
rect 14361 -3081 14373 -3047
rect 12381 -3087 14373 -3081
rect 14439 -3047 16431 -3041
rect 14439 -3081 14451 -3047
rect 16419 -3081 16431 -3047
rect 14439 -3087 16431 -3081
rect 16497 -3047 18489 -3041
rect 16497 -3081 16509 -3047
rect 18477 -3081 18489 -3047
rect 16497 -3087 18489 -3081
rect 18555 -3047 20547 -3041
rect 18555 -3081 18567 -3047
rect 20535 -3081 20547 -3047
rect 18555 -3087 20547 -3081
rect 20613 -3047 22605 -3041
rect 20613 -3081 20625 -3047
rect 22593 -3081 22605 -3047
rect 20613 -3087 22605 -3081
rect 22671 -3047 24663 -3041
rect 22671 -3081 22683 -3047
rect 24651 -3081 24663 -3047
rect 22671 -3087 24663 -3081
rect 24729 -3047 26721 -3041
rect 24729 -3081 24741 -3047
rect 26709 -3081 26721 -3047
rect 24729 -3087 26721 -3081
rect 26787 -3047 28779 -3041
rect 26787 -3081 26799 -3047
rect 28767 -3081 28779 -3047
rect 26787 -3087 28779 -3081
<< properties >>
string FIXED_BBOX -28926 -3166 28926 3166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 30 l 10 m 1 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
