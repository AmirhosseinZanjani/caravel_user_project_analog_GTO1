magic
tech sky130A
magscale 1 2
timestamp 1697806833
<< nwell >>
rect -3254 -4019 3254 4019
<< pmos >>
rect -3058 -3800 -1058 3800
rect -1000 -3800 1000 3800
rect 1058 -3800 3058 3800
<< pdiff >>
rect -3116 3788 -3058 3800
rect -3116 -3788 -3104 3788
rect -3070 -3788 -3058 3788
rect -3116 -3800 -3058 -3788
rect -1058 3788 -1000 3800
rect -1058 -3788 -1046 3788
rect -1012 -3788 -1000 3788
rect -1058 -3800 -1000 -3788
rect 1000 3788 1058 3800
rect 1000 -3788 1012 3788
rect 1046 -3788 1058 3788
rect 1000 -3800 1058 -3788
rect 3058 3788 3116 3800
rect 3058 -3788 3070 3788
rect 3104 -3788 3116 3788
rect 3058 -3800 3116 -3788
<< pdiffc >>
rect -3104 -3788 -3070 3788
rect -1046 -3788 -1012 3788
rect 1012 -3788 1046 3788
rect 3070 -3788 3104 3788
<< nsubdiff >>
rect -3218 3949 -3122 3983
rect 3122 3949 3218 3983
rect -3218 3887 -3184 3949
rect 3184 3887 3218 3949
rect -3218 -3949 -3184 -3887
rect 3184 -3949 3218 -3887
rect -3218 -3983 -3122 -3949
rect 3122 -3983 3218 -3949
<< nsubdiffcont >>
rect -3122 3949 3122 3983
rect -3218 -3887 -3184 3887
rect 3184 -3887 3218 3887
rect -3122 -3983 3122 -3949
<< poly >>
rect -3058 3881 -1058 3897
rect -3058 3847 -3042 3881
rect -1074 3847 -1058 3881
rect -3058 3800 -1058 3847
rect -1000 3881 1000 3897
rect -1000 3847 -984 3881
rect 984 3847 1000 3881
rect -1000 3800 1000 3847
rect 1058 3881 3058 3897
rect 1058 3847 1074 3881
rect 3042 3847 3058 3881
rect 1058 3800 3058 3847
rect -3058 -3847 -1058 -3800
rect -3058 -3881 -3042 -3847
rect -1074 -3881 -1058 -3847
rect -3058 -3897 -1058 -3881
rect -1000 -3847 1000 -3800
rect -1000 -3881 -984 -3847
rect 984 -3881 1000 -3847
rect -1000 -3897 1000 -3881
rect 1058 -3847 3058 -3800
rect 1058 -3881 1074 -3847
rect 3042 -3881 3058 -3847
rect 1058 -3897 3058 -3881
<< polycont >>
rect -3042 3847 -1074 3881
rect -984 3847 984 3881
rect 1074 3847 3042 3881
rect -3042 -3881 -1074 -3847
rect -984 -3881 984 -3847
rect 1074 -3881 3042 -3847
<< locali >>
rect -3218 3949 -3122 3983
rect 3122 3949 3218 3983
rect -3218 3887 -3184 3949
rect 3184 3887 3218 3949
rect -3058 3847 -3042 3881
rect -1074 3847 -1058 3881
rect -1000 3847 -984 3881
rect 984 3847 1000 3881
rect 1058 3847 1074 3881
rect 3042 3847 3058 3881
rect -3104 3788 -3070 3804
rect -3104 -3804 -3070 -3788
rect -1046 3788 -1012 3804
rect -1046 -3804 -1012 -3788
rect 1012 3788 1046 3804
rect 1012 -3804 1046 -3788
rect 3070 3788 3104 3804
rect 3070 -3804 3104 -3788
rect -3058 -3881 -3042 -3847
rect -1074 -3881 -1058 -3847
rect -1000 -3881 -984 -3847
rect 984 -3881 1000 -3847
rect 1058 -3881 1074 -3847
rect 3042 -3881 3058 -3847
rect -3218 -3949 -3184 -3887
rect 3184 -3949 3218 -3887
rect -3218 -3983 -3122 -3949
rect 3122 -3983 3218 -3949
<< viali >>
rect -3042 3847 -1074 3881
rect -984 3847 984 3881
rect 1074 3847 3042 3881
rect -3104 -3788 -3070 3788
rect -1046 -3788 -1012 3788
rect 1012 -3788 1046 3788
rect 3070 -3788 3104 3788
rect -3042 -3881 -1074 -3847
rect -984 -3881 984 -3847
rect 1074 -3881 3042 -3847
<< metal1 >>
rect -3054 3881 -1062 3887
rect -3054 3847 -3042 3881
rect -1074 3847 -1062 3881
rect -3054 3841 -1062 3847
rect -996 3881 996 3887
rect -996 3847 -984 3881
rect 984 3847 996 3881
rect -996 3841 996 3847
rect 1062 3881 3054 3887
rect 1062 3847 1074 3881
rect 3042 3847 3054 3881
rect 1062 3841 3054 3847
rect -3110 3788 -3064 3800
rect -3110 -3788 -3104 3788
rect -3070 -3788 -3064 3788
rect -3110 -3800 -3064 -3788
rect -1052 3788 -1006 3800
rect -1052 -3788 -1046 3788
rect -1012 -3788 -1006 3788
rect -1052 -3800 -1006 -3788
rect 1006 3788 1052 3800
rect 1006 -3788 1012 3788
rect 1046 -3788 1052 3788
rect 1006 -3800 1052 -3788
rect 3064 3788 3110 3800
rect 3064 -3788 3070 3788
rect 3104 -3788 3110 3788
rect 3064 -3800 3110 -3788
rect -3054 -3847 -1062 -3841
rect -3054 -3881 -3042 -3847
rect -1074 -3881 -1062 -3847
rect -3054 -3887 -1062 -3881
rect -996 -3847 996 -3841
rect -996 -3881 -984 -3847
rect 984 -3881 996 -3847
rect -996 -3887 996 -3881
rect 1062 -3847 3054 -3841
rect 1062 -3881 1074 -3847
rect 3042 -3881 3054 -3847
rect 1062 -3887 3054 -3881
<< properties >>
string FIXED_BBOX -3201 -3966 3201 3966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 38 l 10 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
