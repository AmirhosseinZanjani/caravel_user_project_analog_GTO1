magic
tech sky130A
magscale 1 2
timestamp 1694443192
<< error_p >>
rect 229 729 287 735
rect 421 729 479 735
rect 613 729 671 735
rect 805 729 863 735
rect 997 729 1055 735
rect 1189 729 1247 735
rect 1381 729 1439 735
rect 229 695 241 729
rect 421 695 433 729
rect 613 695 625 729
rect 805 695 817 729
rect 997 695 1009 729
rect 1189 695 1201 729
rect 1381 695 1393 729
rect 229 689 287 695
rect 421 689 479 695
rect 613 689 671 695
rect 805 689 863 695
rect 997 689 1055 695
rect 1189 689 1247 695
rect 1381 689 1439 695
rect 133 119 191 125
rect 325 119 383 125
rect 517 119 575 125
rect 709 119 767 125
rect 901 119 959 125
rect 1093 119 1151 125
rect 1285 119 1343 125
rect 133 85 145 119
rect 325 85 337 119
rect 517 85 529 119
rect 709 85 721 119
rect 901 85 913 119
rect 1093 85 1105 119
rect 1285 85 1297 119
rect 133 79 191 85
rect 325 79 383 85
rect 517 79 575 85
rect 709 79 767 85
rect 901 79 959 85
rect 1093 79 1151 85
rect 1285 79 1343 85
use sky130_fd_pr__nfet_01v8_LM9D52  sky130_fd_pr__nfet_01v8_LM9D52_0
timestamp 1694443192
transform 1 0 786 0 1 407
box -839 -460 839 460
<< end >>
