magic
tech sky130A
magscale 1 2
timestamp 1695730805
<< locali >>
rect 1246 -8404 1376 14704
<< metal1 >>
rect 3234 13586 3306 13640
rect 3248 6378 3320 6432
rect 3244 2068 3316 2122
rect 3248 -556 3320 -502
rect 3246 -3180 3318 -3126
rect 3248 -7164 3320 -7110
<< metal4 >>
rect -4844 13668 -4444 13708
rect -4844 13348 -4804 13668
rect -4484 13558 -4444 13668
rect 75 13558 76 13776
rect 1096 13558 1097 13776
rect 3445 13558 3446 13776
rect 4466 13558 4467 13776
rect 8986 13668 9386 13708
rect 8986 13558 9026 13668
rect -4484 13458 1188 13558
rect 3366 13458 9026 13558
rect -4484 13348 -4444 13458
rect -4844 13308 -4444 13348
rect 8986 13348 9026 13458
rect 9346 13348 9386 13668
rect 8986 13308 9386 13348
rect 75 6568 76 6582
rect 1096 6568 1097 6582
rect 3445 6568 3446 6582
rect 4466 6568 4467 6582
rect -4844 6460 -4444 6500
rect -4844 6140 -4804 6460
rect -4484 6350 -4444 6460
rect -2485 6350 -2484 6546
rect -1464 6350 -1463 6546
rect 75 6350 76 6546
rect 1096 6350 1097 6546
rect 1388 6350 1488 6546
rect -4484 6250 1488 6350
rect 3066 6350 3166 6546
rect 3445 6350 3446 6546
rect 4466 6350 4467 6546
rect 6005 6350 6006 6546
rect 7026 6350 7027 6546
rect 8986 6460 9386 6500
rect 8986 6350 9026 6460
rect 3066 6250 9026 6350
rect -4484 6140 -4444 6250
rect -4844 6100 -4444 6140
rect 8986 6140 9026 6250
rect 9346 6140 9386 6460
rect 8986 6100 9386 6140
rect -4844 2360 -4444 2400
rect -4844 2040 -4804 2360
rect -4484 2250 -4444 2360
rect 8986 2360 9386 2400
rect 8986 2250 9026 2360
rect -4484 2150 1188 2250
rect 3366 2150 9026 2250
rect -4484 2040 -4444 2150
rect -4844 2000 -4444 2040
rect 8986 2040 9026 2150
rect 9346 2040 9386 2360
rect 8986 2000 9386 2040
rect -4844 -264 -4444 -224
rect -4844 -584 -4804 -264
rect -4484 -374 -4444 -264
rect 8986 -264 9386 -224
rect 8986 -374 9026 -264
rect -4484 -474 1188 -374
rect 3366 -474 9026 -374
rect -4484 -584 -4444 -474
rect -4844 -624 -4444 -584
rect 75 -662 76 -474
rect 1096 -662 1097 -474
rect 3445 -662 3446 -474
rect 4466 -662 4467 -474
rect 8986 -584 9026 -474
rect 9346 -584 9386 -264
rect 8986 -624 9386 -584
rect -4844 -2888 -4444 -2848
rect -4844 -3208 -4804 -2888
rect -4484 -2998 -4444 -2888
rect 8986 -2888 9386 -2848
rect 8986 -2998 9026 -2888
rect -4484 -3098 1188 -2998
rect 3366 -3098 9026 -2998
rect -4484 -3208 -4444 -3098
rect -4844 -3248 -4444 -3208
rect 75 -3286 76 -3098
rect 1096 -3286 1097 -3098
rect 3445 -3286 3446 -3098
rect 4466 -3286 4467 -3098
rect 8986 -3208 9026 -3098
rect 9346 -3208 9386 -2888
rect 8986 -3248 9386 -3208
rect -4844 -6872 -4444 -6832
rect -4844 -7192 -4804 -6872
rect -4484 -6982 -4444 -6872
rect 8986 -6872 9386 -6832
rect 8986 -6982 9026 -6872
rect -4484 -7082 1188 -6982
rect 3366 -7082 9026 -6982
rect -4484 -7192 -4444 -7082
rect -4844 -7232 -4444 -7192
rect 75 -7270 76 -7082
rect 1096 -7270 1097 -7082
rect 3445 -7270 3446 -7082
rect 4466 -7270 4467 -7082
rect 8986 -7192 9026 -7082
rect 9346 -7192 9386 -6872
rect 8986 -7232 9386 -7192
<< via4 >>
rect -4804 13348 -4484 13668
rect 9026 13348 9346 13668
rect -4804 6140 -4484 6460
rect 9026 6140 9346 6460
rect -4804 2040 -4484 2360
rect 9026 2040 9346 2360
rect -4804 -584 -4484 -264
rect 9026 -584 9346 -264
rect -4804 -3208 -4484 -2888
rect 9026 -3208 9346 -2888
rect -4804 -7192 -4484 -6872
rect 9026 -7192 9346 -6872
<< metal5 >>
rect -4844 13668 -4444 19666
rect -4844 13348 -4804 13668
rect -4484 13348 -4444 13668
rect -4844 6460 -4444 13348
rect -4844 6140 -4804 6460
rect -4484 6140 -4444 6460
rect -4844 2360 -4444 6140
rect -4844 2040 -4804 2360
rect -4484 2040 -4444 2360
rect -4844 -264 -4444 2040
rect -4844 -584 -4804 -264
rect -4484 -584 -4444 -264
rect -4844 -2888 -4444 -584
rect -4844 -3208 -4804 -2888
rect -4484 -3208 -4444 -2888
rect -4844 -6872 -4444 -3208
rect -4844 -7192 -4804 -6872
rect -4484 -7192 -4444 -6872
rect -4844 -9966 -4444 -7192
rect 8986 13668 9386 19666
rect 8986 13348 9026 13668
rect 9346 13348 9386 13668
rect 8986 6460 9386 13348
rect 8986 6140 9026 6460
rect 9346 6140 9386 6460
rect 8986 2360 9386 6140
rect 8986 2040 9026 2360
rect 9346 2040 9386 2360
rect 8986 -264 9386 2040
rect 8986 -584 9026 -264
rect 9346 -584 9386 -264
rect 8986 -2888 9386 -584
rect 8986 -3208 9026 -2888
rect 9346 -3208 9386 -2888
rect 8986 -6872 9386 -3208
rect 8986 -7192 9026 -6872
rect 9346 -7192 9386 -6872
rect 8986 -9966 9386 -7192
use capbank_1  capbank_1_0
timestamp 1695720837
transform 1 0 1288 0 -1 2250
box -1292 0 3258 1624
use capbank_2  capbank_2_0
timestamp 1695721010
transform 1 0 1288 0 -1 -374
box -2572 0 4538 1624
use capbank_4  capbank_4_0
timestamp 1695721417
transform 1 0 1288 0 -1 -2998
box -2572 0 4538 2984
use capbank_8  capbank_8_0
timestamp 1695721793
transform 1 0 1288 0 -1 -6982
box -5132 0 7098 2984
use capbank_16  capbank_16_0
timestamp 1695726168
transform 1 0 1288 0 1 13458
box -5132 0 7098 6208
use capbank_16  capbank_16_1
timestamp 1695726168
transform 1 0 1288 0 1 6250
box -5132 0 7098 6208
<< labels >>
flabel metal5 8986 13668 9386 19666 0 FreeSans 1600 90 0 0 vp_cap
port 1 nsew
flabel metal5 -4844 13668 -4444 19666 0 FreeSans 1600 90 0 0 vn_cap
port 2 nsew
flabel metal1 3244 2068 3316 2122 0 FreeSans 160 0 0 0 tune[0]
port 3 nsew
flabel metal1 3248 -556 3320 -502 0 FreeSans 160 0 0 0 tune[1]
port 4 nsew
flabel metal1 3246 -3180 3318 -3126 0 FreeSans 160 0 0 0 tune[2]
port 5 nsew
flabel metal1 3248 -7164 3320 -7110 0 FreeSans 160 0 0 0 tune[3]
port 6 nsew
flabel metal1 3248 6378 3320 6432 0 FreeSans 160 0 0 0 tune[4]
port 7 nsew
flabel metal1 3234 13586 3306 13640 0 FreeSans 160 0 0 0 tune[5]
port 8 nsew
flabel locali 1246 -8404 1376 14704 0 FreeSans 160 0 0 0 vss_cap
port 0 nsew
<< end >>
