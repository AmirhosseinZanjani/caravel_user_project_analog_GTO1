magic
tech sky130A
magscale 1 2
timestamp 1699606472
<< pwell >>
rect -54 4297 66178 4874
rect -18 -16 52 30
<< locali >>
rect 15968 20364 49776 20368
rect 15968 20200 50350 20364
rect 15958 19986 50350 20200
rect 15958 19982 40076 19986
rect 15958 19934 25410 19982
rect 15958 19810 17684 19934
rect 25364 19900 25410 19934
rect 25852 19934 40076 19982
rect 25852 19900 25908 19934
rect 25364 19896 25908 19900
rect 40040 19904 40076 19934
rect 40518 19934 50350 19986
rect 40518 19904 40536 19934
rect 40040 19890 40536 19904
rect 15958 19808 16642 19810
rect 18680 19808 22714 19850
rect 22796 19808 33008 19850
rect 33086 19808 43300 19850
rect 43376 19808 47404 19850
rect 48410 19808 50350 19934
rect 15958 19290 16598 19808
rect 15958 13226 16482 19290
rect 49488 19284 50350 19808
rect 49606 13234 50350 19284
rect 15958 12714 16594 13226
rect 49492 12716 50350 13234
rect 15958 12706 16638 12714
rect 17300 12706 17732 12714
rect 15958 12640 17732 12706
rect 48356 12640 50350 12716
rect 15956 11970 50354 12640
rect -54 4322 66178 4874
rect -54 4276 -8 4322
rect 62 4318 66178 4322
rect 62 4297 66010 4318
rect -54 2772 10 4276
rect 696 4190 1558 4297
rect 2217 4195 10360 4236
rect 16623 4195 22712 4234
rect 26913 4195 30934 4240
rect 35145 4195 39170 4234
rect 43361 4195 49462 4230
rect 64604 4194 65466 4297
rect 66086 4297 66178 4318
rect 66086 4246 66170 4297
rect -54 1990 138 2772
rect 66064 2748 66170 4246
rect -54 54 10 1990
rect 65940 1966 66170 2748
rect -54 38 84 54
rect -54 -8 -4 38
rect 66 18 84 38
rect 692 18 1554 122
rect 13140 18 13654 116
rect 15308 18 15822 114
rect 23378 18 23702 118
rect 25638 18 25962 116
rect 33000 22 33108 24
rect 33000 18 33018 22
rect 66 10 24782 18
rect 66 -8 14486 10
rect -54 -26 14486 -8
rect 14554 -18 24782 10
rect 24850 -16 33018 18
rect 33070 18 33108 22
rect 39966 18 40290 118
rect 42056 18 42380 116
rect 50242 18 50684 120
rect 51526 24 51610 38
rect 51526 18 51538 24
rect 33070 16 51538 18
rect 33070 -16 41236 16
rect 24850 -18 41236 -16
rect 14554 -26 41236 -18
rect -54 -44 41236 -26
rect 41310 -16 51538 16
rect 51592 18 51610 24
rect 52220 18 52662 120
rect 64578 18 65440 120
rect 66064 54 66170 1966
rect 66026 36 66170 54
rect 66026 18 66036 36
rect 51592 -14 66036 18
rect 66094 18 66170 36
rect 66094 -14 66172 18
rect 51592 -16 66172 -14
rect 41310 -44 66172 -16
rect -54 -114 66172 -44
rect -66 -122 66170 -114
rect -66 -296 66168 -122
<< viali >>
rect 25410 19900 25852 19982
rect 40076 19904 40518 19986
rect -8 4276 62 4322
rect 66010 4246 66086 4318
rect -4 -8 66 38
rect 14486 -26 14554 10
rect 24782 -18 24850 18
rect 33018 -16 33070 22
rect 41236 -44 41310 16
rect 51538 -16 51592 24
rect 66036 -14 66094 36
<< metal1 >>
rect 19376 22514 46358 23186
rect 19376 19802 19706 22514
rect 23654 21478 42456 21872
rect 23650 21474 42456 21478
rect 23650 19798 24006 21474
rect 42088 21192 42456 21474
rect 27604 20340 38328 20726
rect 25400 19884 25410 20020
rect 25858 19884 25868 20020
rect 27606 19790 27912 20340
rect 29642 19754 29652 19848
rect 30000 19754 30010 19848
rect 35748 19742 35758 19836
rect 36106 19742 36116 19836
rect 37988 19806 38326 20340
rect 40058 19892 40068 20048
rect 40516 19986 40526 20048
rect 40518 19904 40526 19986
rect 40516 19892 40526 19904
rect 42118 19792 42456 21192
rect 45996 19796 46326 22514
rect 24736 16082 24746 16434
rect 24864 16082 24874 16434
rect 28866 16062 28876 16414
rect 28994 16062 29004 16414
rect 32956 16068 32966 16420
rect 33084 16068 33094 16420
rect 37088 16052 37098 16404
rect 37216 16052 37226 16404
rect 41200 16044 41210 16396
rect 41328 16044 41338 16396
rect 18592 13956 18602 14204
rect 18666 13956 18676 14204
rect 22704 13960 22714 14208
rect 22778 13960 22788 14208
rect 26812 13950 26822 14198
rect 26886 13950 26896 14198
rect 30924 13952 30934 14200
rect 30998 13952 31008 14200
rect 35056 13960 35066 14208
rect 35130 13960 35140 14208
rect 39162 13970 39172 14218
rect 39236 13970 39246 14218
rect 43290 13970 43300 14218
rect 43364 13970 43374 14218
rect 47394 13946 47404 14194
rect 47468 13946 47478 14194
rect 45356 13172 45366 13290
rect 45418 13172 45428 13290
rect 20660 12998 20670 13116
rect 20722 12998 20732 13116
rect 29704 12718 29714 12776
rect 26912 12716 29714 12718
rect 18680 12680 22714 12716
rect 22796 12682 29714 12716
rect 30062 12718 30072 12776
rect 35792 12718 35802 12772
rect 30062 12682 35802 12718
rect 22796 12680 35802 12682
rect 21670 12294 21998 12680
rect 21670 11396 22002 12294
rect 25610 12192 25942 12680
rect 35792 12678 35802 12680
rect 36150 12718 36160 12772
rect 36150 12680 37122 12718
rect 36150 12678 36160 12680
rect 40072 12192 40372 12728
rect 43376 12680 47400 12718
rect 25610 11920 40388 12192
rect 40072 11916 40372 11920
rect 44204 11396 44586 12680
rect 21670 11354 44586 11396
rect 21674 11096 44586 11354
rect 4896 7786 61096 8520
rect 4906 4790 5322 7786
rect 9100 6396 57056 7008
rect 9104 5292 9524 6396
rect 11134 5698 54772 5702
rect -20 4322 2130 4328
rect -20 4276 -8 4322
rect 62 4276 2130 4322
rect -20 4188 2130 4276
rect 4906 4174 5326 4790
rect 9104 4186 9526 5292
rect 11134 5034 54896 5698
rect 11146 4160 11584 5034
rect 12404 3892 12414 4100
rect 12514 3892 12524 4100
rect 16530 4052 16540 4158
rect 16624 4052 16634 4158
rect 17432 4124 17442 4234
rect 17798 4124 17808 4234
rect 21496 4132 21506 4242
rect 21862 4132 21872 4242
rect 29722 4154 29732 4236
rect 29898 4154 29908 4236
rect 31698 4186 31708 4268
rect 31942 4186 31952 4268
rect 33610 4200 33620 4282
rect 33854 4200 33864 4282
rect 35958 4158 35968 4240
rect 36134 4158 36144 4240
rect 44098 4130 44108 4240
rect 44464 4130 44474 4240
rect 48194 4122 48204 4232
rect 48560 4122 48570 4232
rect 54454 4190 54896 5034
rect 56614 4174 57056 6396
rect 60588 4192 61096 7786
rect 63957 4318 66102 4334
rect 63957 4246 66010 4318
rect 66086 4246 66102 4318
rect 63957 4195 66102 4246
rect 49456 3974 49466 4086
rect 49554 3974 49564 4086
rect 53572 3978 53582 4090
rect 53670 3978 53680 4090
rect 78 2350 88 2448
rect 160 2350 170 2448
rect 4176 2348 4186 2446
rect 4258 2348 4268 2446
rect 8298 2358 8308 2456
rect 8380 2358 8390 2456
rect 57696 2350 57706 2448
rect 57778 2350 57788 2448
rect 61828 2352 61838 2450
rect 61910 2352 61920 2450
rect 65920 2332 65930 2430
rect 66002 2332 66012 2430
rect 22712 1782 22722 1880
rect 22794 1782 22804 1880
rect 28884 1736 28894 1834
rect 28966 1736 28976 1834
rect 37122 1736 37132 1834
rect 37204 1736 37214 1834
rect 43292 1760 43302 1858
rect 43374 1760 43384 1858
rect 16538 1042 16548 1140
rect 16620 1042 16630 1140
rect 20646 1042 20656 1140
rect 20728 1042 20738 1140
rect 26822 988 26832 1086
rect 26904 988 26914 1086
rect 30948 966 30958 1064
rect 31030 966 31040 1064
rect 35060 950 35070 1048
rect 35142 950 35152 1048
rect 39158 958 39168 1056
rect 39240 958 39250 1056
rect 45358 974 45368 1072
rect 45440 974 45450 1072
rect 49450 968 49460 1066
rect 49532 968 49542 1066
rect 2132 284 2142 382
rect 2214 284 2224 382
rect 6250 290 6260 388
rect 6332 290 6342 388
rect 10356 292 10366 390
rect 10438 292 10448 390
rect 18600 352 18610 450
rect 18682 352 18692 450
rect 22710 348 22720 446
rect 22792 348 22802 446
rect 43300 348 43310 446
rect 43382 348 43392 446
rect 47404 348 47414 446
rect 47486 348 47496 446
rect 55634 430 55644 528
rect 55716 430 55726 528
rect 59748 430 59758 528
rect 59830 430 59840 528
rect 63854 418 63864 516
rect 63936 418 63946 516
rect 14478 176 14488 274
rect 14560 176 14570 274
rect 24776 198 24786 296
rect 24858 198 24868 296
rect 33004 178 33014 236
rect 33070 178 33080 236
rect 41222 172 41232 286
rect 41314 172 41324 286
rect 51528 170 51538 226
rect 51592 170 51602 226
rect -18 38 2144 122
rect 2858 118 3278 144
rect 6866 134 7286 150
rect 6864 118 7296 134
rect 2201 85 4888 118
rect 5794 85 9008 118
rect 9672 85 10375 118
rect 11150 116 11570 120
rect -18 -8 -4 38
rect 66 -8 2144 38
rect -18 -20 2144 -8
rect 2858 -282 3278 85
rect 2858 -4564 3280 -282
rect 6864 -674 7296 85
rect 6860 -2684 7296 -674
rect 11140 -728 11576 116
rect 16623 85 22702 118
rect 26896 84 30948 116
rect 35145 85 39178 120
rect 43377 85 49470 118
rect 54336 116 54772 128
rect 14478 10 14488 38
rect 14478 -26 14486 10
rect 14478 -60 14488 -26
rect 14560 -60 14570 38
rect 24772 -60 24782 38
rect 24854 -60 24864 38
rect 33006 -28 33016 30
rect 33072 -28 33082 30
rect 41220 -56 41230 30
rect 41312 -56 41322 30
rect 51526 -18 51538 38
rect 51592 -18 51610 38
rect 51526 -38 51610 -18
rect 11140 -1288 11578 -728
rect 54336 -1288 54790 116
rect 11140 -1804 54790 -1288
rect 58632 -2684 59060 128
rect 6860 -3222 59060 -2684
rect 6860 -3236 58954 -3222
rect 62760 -4564 63178 140
rect 63960 36 66102 124
rect 63960 -14 66036 36
rect 66094 -14 66102 36
rect 63960 -26 66102 -14
rect 2858 -5182 63178 -4564
rect 2858 -5190 63158 -5182
<< via1 >>
rect 25410 19982 25858 20020
rect 25410 19900 25852 19982
rect 25852 19900 25858 19982
rect 25410 19884 25858 19900
rect 29652 19754 30000 19848
rect 35758 19742 36106 19836
rect 40068 19986 40516 20048
rect 40068 19904 40076 19986
rect 40076 19904 40516 19986
rect 40068 19892 40516 19904
rect 24746 16082 24864 16434
rect 28876 16062 28994 16414
rect 32966 16068 33084 16420
rect 37098 16052 37216 16404
rect 41210 16044 41328 16396
rect 18602 13956 18666 14204
rect 22714 13960 22778 14208
rect 26822 13950 26886 14198
rect 30934 13952 30998 14200
rect 35066 13960 35130 14208
rect 39172 13970 39236 14218
rect 43300 13970 43364 14218
rect 47404 13946 47468 14194
rect 45366 13172 45418 13290
rect 20670 12998 20722 13116
rect 29714 12682 30062 12776
rect 35802 12678 36150 12772
rect 12414 3892 12514 4100
rect 16540 4052 16624 4158
rect 17442 4124 17798 4234
rect 21506 4132 21862 4242
rect 29732 4154 29898 4236
rect 31708 4186 31942 4268
rect 33620 4200 33854 4282
rect 35968 4158 36134 4240
rect 44108 4130 44464 4240
rect 48204 4122 48560 4232
rect 49466 3974 49554 4086
rect 53582 3978 53670 4090
rect 88 2350 160 2448
rect 4186 2348 4258 2446
rect 8308 2358 8380 2456
rect 57706 2350 57778 2448
rect 61838 2352 61910 2450
rect 65930 2332 66002 2430
rect 22722 1782 22794 1880
rect 28894 1736 28966 1834
rect 37132 1736 37204 1834
rect 43302 1760 43374 1858
rect 16548 1042 16620 1140
rect 20656 1042 20728 1140
rect 26832 988 26904 1086
rect 30958 966 31030 1064
rect 35070 950 35142 1048
rect 39168 958 39240 1056
rect 45368 974 45440 1072
rect 49460 968 49532 1066
rect 2142 284 2214 382
rect 6260 290 6332 388
rect 10366 292 10438 390
rect 18610 352 18682 450
rect 22720 348 22792 446
rect 43310 348 43382 446
rect 47414 348 47486 446
rect 55644 430 55716 528
rect 59758 430 59830 528
rect 63864 418 63936 516
rect 14488 176 14560 274
rect 24786 198 24858 296
rect 33014 178 33070 236
rect 41232 172 41314 286
rect 51538 170 51592 226
rect 14488 10 14560 38
rect 14488 -26 14554 10
rect 14554 -26 14560 10
rect 14488 -60 14560 -26
rect 24782 18 24854 38
rect 24782 -18 24850 18
rect 24850 -18 24854 18
rect 24782 -60 24854 -18
rect 33016 22 33072 30
rect 33016 -16 33018 22
rect 33018 -16 33070 22
rect 33070 -16 33072 22
rect 33016 -28 33072 -16
rect 41230 16 41312 30
rect 41230 -44 41236 16
rect 41236 -44 41310 16
rect 41310 -44 41312 16
rect 41230 -56 41312 -44
rect 51538 24 51592 38
rect 51538 -16 51592 24
rect 51538 -18 51592 -16
<< metal2 >>
rect 40068 20048 40516 20058
rect 25410 20020 25858 20030
rect 25858 19884 25860 19944
rect 25410 19874 25860 19884
rect 40068 19882 40516 19892
rect 25412 16634 25860 19874
rect 29652 19848 30000 19858
rect 29648 19754 29652 19772
rect 35758 19836 36106 19846
rect 30000 19754 30004 19772
rect 29648 19284 30004 19754
rect 35754 19742 35758 19744
rect 36106 19742 36110 19744
rect 35754 19284 36110 19742
rect 29648 18990 36110 19284
rect 29648 18986 35736 18990
rect 40072 16634 40516 19882
rect 24738 16434 41378 16634
rect 24738 16082 24746 16434
rect 24864 16420 41378 16434
rect 24864 16414 32966 16420
rect 24864 16082 28876 16414
rect 24738 16062 28876 16082
rect 28994 16068 32966 16414
rect 33084 16404 41378 16420
rect 33084 16068 37098 16404
rect 28994 16062 37098 16068
rect 24738 16052 37098 16062
rect 37216 16396 41378 16404
rect 37216 16052 41210 16396
rect 24738 16044 41210 16052
rect 41328 16044 41378 16396
rect 24738 15988 41378 16044
rect 40072 15984 40516 15988
rect 18596 14208 31054 14268
rect 18596 14204 22714 14208
rect 18596 13956 18602 14204
rect 18666 13960 22714 14204
rect 22778 14200 31054 14208
rect 22778 14198 30934 14200
rect 22778 13960 26822 14198
rect 18666 13956 26822 13960
rect 18596 13950 26822 13956
rect 26886 13952 30934 14198
rect 30998 13952 31054 14200
rect 26886 13950 31054 13952
rect 18596 13876 31054 13950
rect 35046 14218 47508 14234
rect 35046 14208 39172 14218
rect 35046 13960 35066 14208
rect 35130 13970 39172 14208
rect 39236 13970 43300 14218
rect 43364 14194 47508 14218
rect 43364 13970 47404 14194
rect 35130 13960 47404 13970
rect 35046 13946 47404 13960
rect 47468 13946 47508 14194
rect 35046 13884 47508 13946
rect 12410 10666 12828 10676
rect 12410 10282 12828 10292
rect 12414 4110 12512 10282
rect 16540 9078 16620 9090
rect 18616 9078 18662 13876
rect 45368 13300 45426 13326
rect 45366 13290 45426 13300
rect 20670 13116 20722 13126
rect 20670 12988 20722 12998
rect 19748 10662 20166 10672
rect 20676 10638 20712 12988
rect 29714 12974 36160 13272
rect 45418 13172 45426 13290
rect 45366 13162 45426 13172
rect 29714 12776 30070 12974
rect 35804 12782 36160 12974
rect 30062 12682 30070 12776
rect 35802 12776 36160 12782
rect 35802 12772 36150 12776
rect 29714 12672 30062 12682
rect 35802 12668 36150 12678
rect 20166 10290 32068 10638
rect 33556 10636 33992 10650
rect 45368 10644 45426 13162
rect 44996 10636 45426 10644
rect 33556 10634 45458 10636
rect 19748 10278 20166 10288
rect 16540 8766 18666 9078
rect 16540 4520 16620 8766
rect 18616 8762 18662 8766
rect 31630 6730 32018 10290
rect 33556 10288 44996 10634
rect 16540 4168 16622 4520
rect 31630 4268 32040 6730
rect 17442 4234 17798 4244
rect 16540 4158 16624 4168
rect 12414 4100 12514 4110
rect 16540 4042 16624 4052
rect 21506 4242 21862 4252
rect 17798 4124 17800 4206
rect 12414 3882 12514 3892
rect 17442 3770 17800 4124
rect 21502 4132 21506 4210
rect 21502 4122 21862 4132
rect 29652 4236 29964 4246
rect 29652 4154 29732 4236
rect 29898 4154 29964 4236
rect 21502 3770 21860 4122
rect 29652 3784 29964 4154
rect 31630 4186 31708 4268
rect 31942 4186 32040 4268
rect 31630 4140 32040 4186
rect 33556 4282 33992 10288
rect 45414 10288 45458 10634
rect 44996 10250 45414 10260
rect 47432 9100 47470 13884
rect 53592 10644 53696 10652
rect 53260 10634 53696 10644
rect 53678 10260 53696 10634
rect 53260 10250 53696 10260
rect 47424 8788 49550 9100
rect 47432 8762 47470 8788
rect 33556 4200 33620 4282
rect 33854 4200 33966 4282
rect 33556 4146 33966 4200
rect 35908 4240 36232 4250
rect 35908 4158 35968 4240
rect 36134 4158 36232 4240
rect 35908 3784 36232 4158
rect 44108 4240 44464 4250
rect 44108 4120 44464 4130
rect 48204 4232 48560 4242
rect 17442 3526 21866 3770
rect 29652 3578 36232 3784
rect 35908 3572 36232 3578
rect 44104 3706 44416 4120
rect 48204 4112 48560 4122
rect 48212 3706 48524 4112
rect 49468 4096 49548 8788
rect 53592 4100 53696 10250
rect 49466 4086 49554 4096
rect 49466 3964 49554 3974
rect 53582 4090 53696 4100
rect 53670 3978 53672 4090
rect 53582 3972 53672 3978
rect 53582 3968 53670 3972
rect 44104 3544 48524 3706
rect 88 2456 8382 2500
rect 57708 2458 65980 2478
rect 88 2448 8308 2456
rect 160 2446 8308 2448
rect 160 2350 4186 2446
rect 88 2340 160 2350
rect 4258 2358 8308 2446
rect 8380 2358 8382 2456
rect 4258 2350 8382 2358
rect 57706 2450 65980 2458
rect 57706 2448 61838 2450
rect 57778 2352 61838 2448
rect 61910 2440 65980 2450
rect 61910 2430 66002 2440
rect 61910 2352 65930 2430
rect 57778 2350 65930 2352
rect 8308 2348 8380 2350
rect 4186 2338 4258 2348
rect 57706 2340 65930 2350
rect 57708 2332 65930 2340
rect 57708 2322 66002 2332
rect 57708 2312 65980 2322
rect 22722 1880 43436 1924
rect 22794 1858 43436 1880
rect 22794 1834 43302 1858
rect 22794 1782 28894 1834
rect 22722 1736 28894 1782
rect 28966 1736 37132 1834
rect 37204 1760 43302 1834
rect 43374 1760 43436 1858
rect 37204 1736 43436 1760
rect 22722 1688 43436 1736
rect 16548 1140 16620 1150
rect 20656 1140 20728 1150
rect 16620 1042 20656 1138
rect 16548 1032 16620 1042
rect 20656 1032 20728 1042
rect 26780 1086 39308 1144
rect 26780 988 26832 1086
rect 26904 1064 39308 1086
rect 26904 988 30958 1064
rect 26780 966 30958 988
rect 31030 1056 39308 1064
rect 31030 1048 39168 1056
rect 31030 966 35070 1048
rect 26780 950 35070 966
rect 35142 958 39168 1048
rect 39240 958 39308 1056
rect 45362 1076 49520 1090
rect 45362 1072 49532 1076
rect 45362 980 45368 1072
rect 45440 1066 49532 1072
rect 45440 980 49460 1066
rect 45368 964 45440 974
rect 49460 958 49532 968
rect 35142 950 39308 958
rect 26780 916 39308 950
rect 55644 534 55716 538
rect 59758 534 59830 538
rect 55644 528 63948 534
rect 18610 450 22792 464
rect 2142 388 2214 392
rect 6260 388 6332 398
rect 10366 390 10438 400
rect 2142 382 6260 388
rect 2214 290 6260 382
rect 6332 292 10366 388
rect 10438 292 10468 388
rect 18682 446 22792 450
rect 18682 352 22720 446
rect 18610 342 18682 352
rect 43310 446 43382 456
rect 22720 338 22792 348
rect 43296 348 43310 436
rect 47414 446 47486 456
rect 43382 348 47414 436
rect 55716 430 59758 528
rect 59830 516 63948 528
rect 59830 430 63864 516
rect 55644 420 55716 430
rect 59758 420 59830 430
rect 63936 430 63948 516
rect 63864 408 63936 418
rect 43296 338 47486 348
rect 43296 324 47478 338
rect 6332 290 10468 292
rect 2214 284 10468 290
rect 24786 296 24858 306
rect 2142 274 2214 284
rect 6260 280 6332 284
rect 10366 282 10438 284
rect 14488 274 14560 284
rect 14488 166 14560 176
rect 24782 198 24786 288
rect 41232 286 41314 296
rect 33022 246 33062 250
rect 24782 188 24858 198
rect 33014 236 33070 246
rect 14488 48 14558 166
rect 14488 38 14560 48
rect 14488 -70 14560 -60
rect 24782 38 24856 188
rect 33014 168 33070 178
rect 51548 236 51582 266
rect 33022 40 33062 168
rect 41232 40 41314 172
rect 51538 226 51592 236
rect 51538 160 51592 170
rect 51548 48 51582 160
rect 24854 -60 24856 38
rect 33016 30 33072 40
rect 33016 -38 33072 -28
rect 41230 30 41314 40
rect 41312 -20 41314 30
rect 51538 38 51592 48
rect 51538 -28 51592 -18
rect 24782 -70 24854 -60
rect 41230 -66 41312 -56
<< via2 >>
rect 12410 10292 12828 10666
rect 19748 10288 20166 10662
rect 44996 10260 45414 10634
rect 53260 10260 53678 10634
<< metal3 >>
rect 53318 13868 54288 13872
rect 53260 13844 54288 13868
rect 12048 13798 12840 13800
rect 11810 13348 11820 13798
rect 12362 13348 12874 13798
rect 53260 13394 53742 13844
rect 54284 13394 54294 13844
rect 53260 13376 54288 13394
rect 12410 10671 12832 13348
rect 12400 10666 12838 10671
rect 12400 10292 12410 10666
rect 12828 10656 12838 10666
rect 16318 10656 16328 11780
rect 12828 10292 16328 10656
rect 12400 10287 12838 10292
rect 16318 10258 16328 10292
rect 17376 10656 17386 11780
rect 19738 10662 20176 10667
rect 19738 10656 19748 10662
rect 17376 10292 19748 10656
rect 17376 10258 17386 10292
rect 19738 10288 19748 10292
rect 20166 10288 20176 10662
rect 48684 10652 48694 11682
rect 19738 10283 20176 10288
rect 44958 10634 48694 10652
rect 44958 10260 44996 10634
rect 45414 10260 48694 10634
rect 44958 10242 48694 10260
rect 48684 10160 48694 10242
rect 49742 10652 49752 11682
rect 53260 10652 53718 13376
rect 49742 10634 53718 10652
rect 49742 10260 53260 10634
rect 53678 10260 53718 10634
rect 49742 10255 53688 10260
rect 49742 10242 53686 10255
rect 49742 10160 49752 10242
<< via3 >>
rect 11820 13348 12362 13798
rect 53742 13394 54284 13844
rect 16328 10258 17376 11780
rect 48694 10160 49742 11682
<< metal4 >>
rect 4722 13799 12348 18118
rect 16306 15638 17432 15654
rect 16306 15454 52992 15638
rect 16306 14780 51678 15454
rect 52972 14780 52992 15454
rect 16306 14656 52992 14780
rect 4722 13798 12363 13799
rect 4722 13370 11820 13798
rect 11819 13348 11820 13370
rect 12362 13348 12363 13798
rect 11819 13347 12363 13348
rect 16306 11780 17432 14656
rect 53752 13845 61378 18130
rect 53741 13844 61378 13845
rect 53741 13394 53742 13844
rect 54284 13394 61378 13844
rect 53741 13393 61378 13394
rect 53752 13382 61378 13393
rect 16306 10258 16328 11780
rect 17376 10258 17432 11780
rect 16306 10218 17432 10258
rect 48693 11682 49743 11683
rect 48693 10160 48694 11682
rect 49742 10160 49743 11682
rect 48693 10159 49743 10160
<< via4 >>
rect 51678 14780 52972 15454
rect 48694 10160 49742 11682
<< mimcap2 >>
rect 5446 15388 11812 17310
rect 5446 14714 10340 15388
rect 11634 14714 11812 15388
rect 5446 14386 11812 14714
rect 54476 15434 60842 17322
rect 54476 14760 54588 15434
rect 55882 14760 60842 15434
rect 54476 14398 60842 14760
<< mimcap2contact >>
rect 10340 14714 11634 15388
rect 54588 14760 55882 15434
<< metal5 >>
rect 10124 15388 49806 15628
rect 10124 14714 10340 15388
rect 11634 14714 49806 15388
rect 10124 14648 49806 14714
rect 51454 15620 55114 15638
rect 51454 15454 56160 15620
rect 51454 14780 51678 15454
rect 52972 15434 56160 15454
rect 52972 14780 54588 15434
rect 51454 14760 54588 14780
rect 55882 14760 56160 15434
rect 51454 14668 56160 14760
rect 52500 14650 56160 14668
rect 48694 11706 49770 14648
rect 48670 11682 49770 11706
rect 48670 10160 48694 11682
rect 49742 10160 49770 11682
rect 48670 10136 49766 10160
use sky130_fd_pr__nfet_01v8_NJ4FLX#0  sky130_fd_pr__nfet_01v8_NJ4FLX_0
timestamp 1699485026
transform 1 0 33042 0 1 2157
box -33095 -2210 33095 2210
use sky130_fd_pr__pfet_01v8_T2K7LE#0  sky130_fd_pr__pfet_01v8_T2K7LE_0
timestamp 1699523894
transform 1 0 33041 0 1 16261
box -16631 -3719 16631 3719
<< labels >>
rlabel metal2 21594 388 21594 388 1 Tail1
rlabel metal2 17154 8874 17154 8874 1 NodeB
rlabel metal2 48026 8942 48026 8942 1 NodeA
rlabel metal2 33698 3704 33698 3704 1 BiasTail
port 10 n
rlabel metal1 17842 -1590 17842 -1590 1 BiasN2
port 9 n
rlabel locali 182 4734 182 4734 1 vss
port 8 n
rlabel metal1 3904 -5042 3904 -5042 1 BiasN1
port 7 n
rlabel metal3 46640 10438 46640 10438 1 ON
port 6 n
rlabel metal3 14012 10468 14012 10468 1 OP
port 5 n
rlabel metal1 24922 22916 24922 22916 1 BiasP1
port 2 n
rlabel metal1 28280 21630 28280 21630 1 BiasP2
port 1 n
rlabel metal2 46574 3618 46574 3618 1 InN
port 4 n
rlabel metal2 19616 3654 19616 3654 1 InP
port 3 n
rlabel locali 17184 20244 17184 20244 1 vdd
port 0 n
<< end >>
